////////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   / 
// /___/  \  /    Vendor: Xilinx 
// \   \   \/     Version : 1.8
//  \   \         Application : Virtex-6 FPGA GTX Transceiver Wizard 
//  /   /         Filename : snap12_t20r20_top.v
// /___/   /\     Timestamp : 
// \   \  /  \ 
//  \___\/\___\ 
//
//
// Module SNAP12_T20R20_TOP
// Generated by Xilinx Virtex-6 FPGA GTX Transceiver Wizard
// 

`timescale 1ns / 1ps
`define DLY #1


//***********************************Entity Declaration************************

module SNAP12_T20R20_TOP #
(
    parameter EXAMPLE_CONFIG_INDEPENDENT_LANES          =   1,   //configuration for frame gen and check
    parameter EXAMPLE_LANE_WITH_START_CHAR              =   0,    // specifies lane with unique start frame char
    parameter EXAMPLE_WORDS_IN_BRAM                     =   512,  // specifies amount of data in BRAM
    parameter EXAMPLE_SIM_GTXRESET_SPEEDUP              =   0,    // simulation setting for GTX SecureIP model
    parameter EXAMPLE_USE_CHIPSCOPE                     =   1,    // Set to 1 to use Chipscope to drive resets
    parameter ALIGNER_WAIT                              =   8'd32 // To set the wait cycles in aligner
)
(
    input wire     ck_160n,
    input wire     ck_160p,
    input wire  [7:0]  RXN,
    input wire  [7:0]  RXP,
    output wire [7:0]  TXN,
    output wire [7:0]  TXP,
    output wire    snap_clk2, ck_160_plllkdet,
    input wire     GTXTXRESET_IN,  // == reset
    input wire     GTXRXRESET_IN,  // == reset
    input   [15:0] SEED_STEP,
    input          gtx_wait,
    input          force_err_wait,
    input   [7:0]  force_err_flag,
    input          snap_commaalign,
    input   [64:0] SEED_BASE,
    output         all_rx_ready, all_tx_ready,
    output  [7:0]  rxdv_snapr, rxcomma_snapr, syncdone_snapt, // my RxDV and Comma
    output  [7:0]  check_ok_snapr, check_bad_snapr, good_byte, bad_byte, lost_byte,
    output [31:0] snap_err0,  // 32-bit wide error count for snap12 tx-rx loop  ___DEFINE THESE IN LOWER LEVELS!
    output [31:0] snap_err1,  // 32-bit wide error count for snap12 tx-rx loop
    output [31:0] snap_err2,  // 32-bit wide error count for snap12 tx-rx loop
    output [31:0] snap_err3,  // 32-bit wide error count for snap12 tx-rx loop
    output [31:0] snap_err4,  // 32-bit wide error count for snap12 tx-rx loop
    output [31:0] snap_err5,  // 32-bit wide error count for snap12 tx-rx loop
    output [31:0] snap_err6,  // 32-bit wide error count for snap12 tx-rx loop
    output [31:0] snap_err7,  // 32-bit wide error count for snap12 tx-rx loop
    output wire [7:0]  rxdv_diff, rxcomma_diff, // diff between my RxDV/Comma and Theirs
    output  [15:0] rxdata_i,
    output  [1:0] RXK_OUT
);


    reg [64:0] seed_in[7:0];
    integer  i;

    initial begin
       for (i = 0; i < 8; i = i + 1) begin
          seed_in[i] = SEED_BASE[64:0] + (((i+1)*2901*SEED_STEP[15:0]) + i << 15);
//	  seed_in[i] = SEED_BASE[64:0];
       end
    end


//************************** Register Declarations ****************************

    reg     [84:0]  ila_in_r;

    reg             gtx0_txresetdone_r;
    reg             gtx0_txresetdone_r2;
// * max_fanout = 1 *
    reg             gtx0_rxresetdone_i_r;
    reg             gtx0_rxresetdone_r;
    reg             gtx0_rxresetdone_r2;
    reg             gtx0_rxresetdone_r3;
    reg             gtx1_txresetdone_r;
    reg             gtx1_txresetdone_r2;
// * max_fanout = 1 *
    reg             gtx1_rxresetdone_i_r;
    reg             gtx1_rxresetdone_r;
    reg             gtx1_rxresetdone_r2;
    reg             gtx1_rxresetdone_r3;
    reg             gtx2_txresetdone_r;
    reg             gtx2_txresetdone_r2;
// * max_fanout = 1 *
    reg             gtx2_rxresetdone_i_r;
    reg             gtx2_rxresetdone_r;
    reg             gtx2_rxresetdone_r2;
    reg             gtx2_rxresetdone_r3;
    reg             gtx3_txresetdone_r;
    reg             gtx3_txresetdone_r2;
// * max_fanout = 1 *
    reg             gtx3_rxresetdone_i_r;
    reg             gtx3_rxresetdone_r;
    reg             gtx3_rxresetdone_r2;
    reg             gtx3_rxresetdone_r3;
    reg             gtx4_txresetdone_r;
    reg             gtx4_txresetdone_r2;
// * max_fanout = 1 *
    reg             gtx4_rxresetdone_i_r;
    reg             gtx4_rxresetdone_r;
    reg             gtx4_rxresetdone_r2;
    reg             gtx4_rxresetdone_r3;
    reg             gtx5_txresetdone_r;
    reg             gtx5_txresetdone_r2;
// * max_fanout = 1 *
    reg             gtx5_rxresetdone_i_r;
    reg             gtx5_rxresetdone_r;
    reg             gtx5_rxresetdone_r2;
    reg             gtx5_rxresetdone_r3;
    reg             gtx6_txresetdone_r;
    reg             gtx6_txresetdone_r2;
// * max_fanout = 1 *
    reg             gtx6_rxresetdone_i_r;
    reg             gtx6_rxresetdone_r;
    reg             gtx6_rxresetdone_r2;
    reg             gtx6_rxresetdone_r3;
    reg             gtx7_txresetdone_r;
    reg             gtx7_txresetdone_r2;
// * max_fanout = 1 *
    reg             gtx7_rxresetdone_i_r;
    reg             gtx7_rxresetdone_r;
    reg             gtx7_rxresetdone_r2;
    reg             gtx7_rxresetdone_r3;
    reg             gtx8_txresetdone_r;
    reg             gtx8_txresetdone_r2;
// * max_fanout = 1 *
    reg             gtx8_rxresetdone_i_r;
    reg             gtx8_rxresetdone_r;
    reg             gtx8_rxresetdone_r2;
    reg             gtx8_rxresetdone_r3;
    reg             gtx9_txresetdone_r;
    reg             gtx9_txresetdone_r2;
// * max_fanout = 1 *
    reg             gtx9_rxresetdone_i_r;
    reg             gtx9_rxresetdone_r;
    reg             gtx9_rxresetdone_r2;
    reg             gtx9_rxresetdone_r3;
    reg             gtx10_txresetdone_r;
    reg             gtx10_txresetdone_r2;
// * max_fanout = 1 *
    reg             gtx10_rxresetdone_i_r;
    reg             gtx10_rxresetdone_r;
    reg             gtx10_rxresetdone_r2;
    reg             gtx10_rxresetdone_r3;
    reg             gtx11_txresetdone_r;
    reg             gtx11_txresetdone_r2;
// * max_fanout = 1 *
    reg             gtx11_rxresetdone_i_r;
    reg             gtx11_rxresetdone_r;
    reg             gtx11_rxresetdone_r2;
    reg             gtx11_rxresetdone_r3;
    //------------------------ MGT Wrapper Wires ------------------------------
    //________________________________________________________________________
    //________________________________________________________________________
    //GTX0   (X0Y0)

    //---------------------- Loopback and Powerdown Ports ----------------------
    wire    [1:0]   gtx0_rxpowerdown_i;
    wire    [1:0]   gtx0_txpowerdown_i;
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire    [1:0]   gtx0_rxchariscomma_i;
    wire    [1:0]   gtx0_rxcharisk_i;
    wire    [1:0]   gtx0_rxdisperr_i;
    wire    [1:0]   gtx0_rxnotintable_i;
    //----------------- Receive Ports - Clock Correction Ports -----------------
    wire    [2:0]   gtx0_rxclkcorcnt_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            gtx0_rxbyterealign_i;
    wire            gtx0_rxcommadet_i;
    wire            gtx0_rxenmcommaalign_i;
    wire            gtx0_rxenpcommaalign_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [15:0]  gtx0_rxdata_i;
    wire            gtx0_rxreset_i;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    wire            gtx0_rxcdrreset_i;
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    wire    [2:0]   gtx0_rxbufstatus_i;
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    wire    [1:0]   gtx0_rxlossofsync_i;
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    wire            gtx0_gtxrxreset_i;
    wire            gtx0_pllrxreset_i;
    wire            gtx0_rxplllkdet_i;
    wire            gtx0_rxresetdone_i;
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    wire            gtx0_rxvalid_i;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    wire            gtx0_rxpolarity_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [15:0]  gtx0_txdata_i;
    wire            gtx0_txoutclk_i;
    wire            gtx0_txreset_i;
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    wire            gtx0_txdlyaligndisable_i;
    wire            gtx0_txdlyalignmonenb_i;
    wire    [7:0]   gtx0_txdlyalignmonitor_i;
    wire            gtx0_txdlyalignreset_i;
    wire            gtx0_txenpmaphasealign_i;
    wire            gtx0_txpmasetphase_i;
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    wire            gtx0_gtxtxreset_i;
    wire            gtx0_txresetdone_i;


    //________________________________________________________________________
    //________________________________________________________________________
    //GTX1   (X0Y1)

    //---------------------- Loopback and Powerdown Ports ----------------------
    wire    [1:0]   gtx1_rxpowerdown_i;
    wire    [1:0]   gtx1_txpowerdown_i;
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire    [1:0]   gtx1_rxchariscomma_i;
    wire    [1:0]   gtx1_rxcharisk_i;
    wire    [1:0]   gtx1_rxdisperr_i;
    wire    [1:0]   gtx1_rxnotintable_i;
    //----------------- Receive Ports - Clock Correction Ports -----------------
    wire    [2:0]   gtx1_rxclkcorcnt_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            gtx1_rxbyterealign_i;
    wire            gtx1_rxcommadet_i;
    wire            gtx1_rxenmcommaalign_i;
    wire            gtx1_rxenpcommaalign_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [15:0]  gtx1_rxdata_i;
    wire            gtx1_rxreset_i;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    wire            gtx1_rxcdrreset_i;
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    wire    [2:0]   gtx1_rxbufstatus_i;
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    wire    [1:0]   gtx1_rxlossofsync_i;
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    wire            gtx1_gtxrxreset_i;
    wire            gtx1_pllrxreset_i;
    wire            gtx1_rxplllkdet_i;
    wire            gtx1_rxresetdone_i;
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    wire            gtx1_rxvalid_i;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    wire            gtx1_rxpolarity_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [15:0]  gtx1_txdata_i;
    wire            gtx1_txoutclk_i;
    wire            gtx1_txreset_i;
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    wire            gtx1_txdlyaligndisable_i;
    wire            gtx1_txdlyalignmonenb_i;
    wire    [7:0]   gtx1_txdlyalignmonitor_i;
    wire            gtx1_txdlyalignreset_i;
    wire            gtx1_txenpmaphasealign_i;
    wire            gtx1_txpmasetphase_i;
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    wire            gtx1_gtxtxreset_i;
    wire            gtx1_txresetdone_i;


    //________________________________________________________________________
    //________________________________________________________________________
    //GTX2   (X0Y2)

    //---------------------- Loopback and Powerdown Ports ----------------------
    wire    [1:0]   gtx2_rxpowerdown_i;
    wire    [1:0]   gtx2_txpowerdown_i;
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire    [1:0]   gtx2_rxchariscomma_i;
    wire    [1:0]   gtx2_rxcharisk_i;
    wire    [1:0]   gtx2_rxdisperr_i;
    wire    [1:0]   gtx2_rxnotintable_i;
    //----------------- Receive Ports - Clock Correction Ports -----------------
    wire    [2:0]   gtx2_rxclkcorcnt_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            gtx2_rxbyterealign_i;
    wire            gtx2_rxcommadet_i;
    wire            gtx2_rxenmcommaalign_i;
    wire            gtx2_rxenpcommaalign_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [15:0]  gtx2_rxdata_i;
    wire            gtx2_rxreset_i;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    wire            gtx2_rxcdrreset_i;
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    wire    [2:0]   gtx2_rxbufstatus_i;
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    wire    [1:0]   gtx2_rxlossofsync_i;
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    wire            gtx2_gtxrxreset_i;
    wire            gtx2_pllrxreset_i;
    wire            gtx2_rxplllkdet_i;
    wire            gtx2_rxresetdone_i;
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    wire            gtx2_rxvalid_i;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    wire            gtx2_rxpolarity_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [15:0]  gtx2_txdata_i;
    wire            gtx2_txoutclk_i;
    wire            gtx2_txreset_i;
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    wire            gtx2_txdlyaligndisable_i;
    wire            gtx2_txdlyalignmonenb_i;
    wire    [7:0]   gtx2_txdlyalignmonitor_i;
    wire            gtx2_txdlyalignreset_i;
    wire            gtx2_txenpmaphasealign_i;
    wire            gtx2_txpmasetphase_i;
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    wire            gtx2_gtxtxreset_i;
    wire            gtx2_txresetdone_i;


    //________________________________________________________________________
    //________________________________________________________________________
    //GTX3   (X0Y3)

    //---------------------- Loopback and Powerdown Ports ----------------------
    wire    [1:0]   gtx3_rxpowerdown_i;
    wire    [1:0]   gtx3_txpowerdown_i;
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire    [1:0]   gtx3_rxchariscomma_i;
    wire    [1:0]   gtx3_rxcharisk_i;
    wire    [1:0]   gtx3_rxdisperr_i;
    wire    [1:0]   gtx3_rxnotintable_i;
    //----------------- Receive Ports - Clock Correction Ports -----------------
    wire    [2:0]   gtx3_rxclkcorcnt_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            gtx3_rxbyterealign_i;
    wire            gtx3_rxcommadet_i;
    wire            gtx3_rxenmcommaalign_i;
    wire            gtx3_rxenpcommaalign_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [15:0]  gtx3_rxdata_i;
    wire            gtx3_rxreset_i;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    wire            gtx3_rxcdrreset_i;
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    wire    [2:0]   gtx3_rxbufstatus_i;
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    wire    [1:0]   gtx3_rxlossofsync_i;
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    wire            gtx3_gtxrxreset_i;
    wire            gtx3_pllrxreset_i;
    wire            gtx3_rxplllkdet_i;
    wire            gtx3_rxresetdone_i;
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    wire            gtx3_rxvalid_i;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    wire            gtx3_rxpolarity_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [15:0]  gtx3_txdata_i;
    wire            gtx3_txoutclk_i;
    wire            gtx3_txreset_i;
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    wire            gtx3_txdlyaligndisable_i;
    wire            gtx3_txdlyalignmonenb_i;
    wire    [7:0]   gtx3_txdlyalignmonitor_i;
    wire            gtx3_txdlyalignreset_i;
    wire            gtx3_txenpmaphasealign_i;
    wire            gtx3_txpmasetphase_i;
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    wire            gtx3_gtxtxreset_i;
    wire            gtx3_txresetdone_i;


    //________________________________________________________________________
    //________________________________________________________________________
    //GTX4   (X0Y4)

    //---------------------- Loopback and Powerdown Ports ----------------------
    wire    [1:0]   gtx4_rxpowerdown_i;
    wire    [1:0]   gtx4_txpowerdown_i;
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire    [1:0]   gtx4_rxchariscomma_i;
    wire    [1:0]   gtx4_rxcharisk_i;
    wire    [1:0]   gtx4_rxdisperr_i;
    wire    [1:0]   gtx4_rxnotintable_i;
    //----------------- Receive Ports - Clock Correction Ports -----------------
    wire    [2:0]   gtx4_rxclkcorcnt_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            gtx4_rxbyterealign_i;
    wire            gtx4_rxcommadet_i;
    wire            gtx4_rxenmcommaalign_i;
    wire            gtx4_rxenpcommaalign_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [15:0]  gtx4_rxdata_i;
    wire            gtx4_rxreset_i;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    wire            gtx4_rxcdrreset_i;
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    wire    [2:0]   gtx4_rxbufstatus_i;
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    wire    [1:0]   gtx4_rxlossofsync_i;
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    wire            gtx4_gtxrxreset_i;
    wire            gtx4_pllrxreset_i;
    wire            gtx4_rxplllkdet_i;
    wire            gtx4_rxresetdone_i;
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    wire            gtx4_rxvalid_i;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    wire            gtx4_rxpolarity_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [15:0]  gtx4_txdata_i;
    wire            gtx4_txoutclk_i;
    wire            gtx4_txreset_i;
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    wire            gtx4_txdlyaligndisable_i;
    wire            gtx4_txdlyalignmonenb_i;
    wire    [7:0]   gtx4_txdlyalignmonitor_i;
    wire            gtx4_txdlyalignreset_i;
    wire            gtx4_txenpmaphasealign_i;
    wire            gtx4_txpmasetphase_i;
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    wire            gtx4_gtxtxreset_i;
    wire            gtx4_txresetdone_i;


    //________________________________________________________________________
    //________________________________________________________________________
    //GTX5   (X0Y5)

    //---------------------- Loopback and Powerdown Ports ----------------------
    wire    [1:0]   gtx5_rxpowerdown_i;
    wire    [1:0]   gtx5_txpowerdown_i;
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire    [1:0]   gtx5_rxchariscomma_i;
    wire    [1:0]   gtx5_rxcharisk_i;
    wire    [1:0]   gtx5_rxdisperr_i;
    wire    [1:0]   gtx5_rxnotintable_i;
    //----------------- Receive Ports - Clock Correction Ports -----------------
    wire    [2:0]   gtx5_rxclkcorcnt_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            gtx5_rxbyterealign_i;
    wire            gtx5_rxcommadet_i;
    wire            gtx5_rxenmcommaalign_i;
    wire            gtx5_rxenpcommaalign_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [15:0]  gtx5_rxdata_i;
    wire            gtx5_rxreset_i;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    wire            gtx5_rxcdrreset_i;
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    wire    [2:0]   gtx5_rxbufstatus_i;
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    wire    [1:0]   gtx5_rxlossofsync_i;
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    wire            gtx5_gtxrxreset_i;
    wire            gtx5_pllrxreset_i;
    wire            gtx5_rxplllkdet_i;
    wire            gtx5_rxresetdone_i;
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    wire            gtx5_rxvalid_i;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    wire            gtx5_rxpolarity_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [15:0]  gtx5_txdata_i;
    wire            gtx5_txoutclk_i;
    wire            gtx5_txreset_i;
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    wire            gtx5_txdlyaligndisable_i;
    wire            gtx5_txdlyalignmonenb_i;
    wire    [7:0]   gtx5_txdlyalignmonitor_i;
    wire            gtx5_txdlyalignreset_i;
    wire            gtx5_txenpmaphasealign_i;
    wire            gtx5_txpmasetphase_i;
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    wire            gtx5_gtxtxreset_i;
    wire            gtx5_txresetdone_i;


    //________________________________________________________________________
    //________________________________________________________________________
    //GTX6   (X0Y6)

    //---------------------- Loopback and Powerdown Ports ----------------------
    wire    [1:0]   gtx6_rxpowerdown_i;
    wire    [1:0]   gtx6_txpowerdown_i;
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire    [1:0]   gtx6_rxchariscomma_i;
    wire    [1:0]   gtx6_rxcharisk_i;
    wire    [1:0]   gtx6_rxdisperr_i;
    wire    [1:0]   gtx6_rxnotintable_i;
    //----------------- Receive Ports - Clock Correction Ports -----------------
    wire    [2:0]   gtx6_rxclkcorcnt_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            gtx6_rxbyterealign_i;
    wire            gtx6_rxcommadet_i;
    wire            gtx6_rxenmcommaalign_i;
    wire            gtx6_rxenpcommaalign_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [15:0]  gtx6_rxdata_i;
    wire            gtx6_rxreset_i;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    wire            gtx6_rxcdrreset_i;
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    wire    [2:0]   gtx6_rxbufstatus_i;
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    wire    [1:0]   gtx6_rxlossofsync_i;
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    wire            gtx6_gtxrxreset_i;
    wire            gtx6_pllrxreset_i;
    wire            gtx6_rxplllkdet_i;
    wire            gtx6_rxresetdone_i;
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    wire            gtx6_rxvalid_i;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    wire            gtx6_rxpolarity_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [15:0]  gtx6_txdata_i;
    wire            gtx6_txoutclk_i;
    wire            gtx6_txreset_i;
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    wire            gtx6_txdlyaligndisable_i;
    wire            gtx6_txdlyalignmonenb_i;
    wire    [7:0]   gtx6_txdlyalignmonitor_i;
    wire            gtx6_txdlyalignreset_i;
    wire            gtx6_txenpmaphasealign_i;
    wire            gtx6_txpmasetphase_i;
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    wire            gtx6_gtxtxreset_i;
    wire            gtx6_txresetdone_i;


    //________________________________________________________________________
    //________________________________________________________________________
    //GTX7   (X0Y7)

    //---------------------- Loopback and Powerdown Ports ----------------------
    wire    [1:0]   gtx7_rxpowerdown_i;
    wire    [1:0]   gtx7_txpowerdown_i;
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire    [1:0]   gtx7_rxchariscomma_i;
    wire    [1:0]   gtx7_rxcharisk_i;
    wire    [1:0]   gtx7_rxdisperr_i;
    wire    [1:0]   gtx7_rxnotintable_i;
    //----------------- Receive Ports - Clock Correction Ports -----------------
    wire    [2:0]   gtx7_rxclkcorcnt_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            gtx7_rxbyterealign_i;
    wire            gtx7_rxcommadet_i;
    wire            gtx7_rxenmcommaalign_i;
    wire            gtx7_rxenpcommaalign_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [15:0]  gtx7_rxdata_i;
    wire            gtx7_rxreset_i;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    wire            gtx7_rxcdrreset_i;
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    wire    [2:0]   gtx7_rxbufstatus_i;
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    wire    [1:0]   gtx7_rxlossofsync_i;
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    wire            gtx7_gtxrxreset_i;
    wire            gtx7_pllrxreset_i;
    wire            gtx7_rxplllkdet_i;
    wire            gtx7_rxresetdone_i;
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    wire            gtx7_rxvalid_i;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    wire            gtx7_rxpolarity_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [15:0]  gtx7_txdata_i;
    wire            gtx7_txoutclk_i;
    wire            gtx7_txreset_i;
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    wire            gtx7_txdlyaligndisable_i;
    wire            gtx7_txdlyalignmonenb_i;
    wire    [7:0]   gtx7_txdlyalignmonitor_i;
    wire            gtx7_txdlyalignreset_i;
    wire            gtx7_txenpmaphasealign_i;
    wire            gtx7_txpmasetphase_i;
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    wire            gtx7_gtxtxreset_i;
    wire            gtx7_txresetdone_i;


    //________________________________________________________________________
    //________________________________________________________________________
    //GTX8   (X0Y8)

    //---------------------- Loopback and Powerdown Ports ----------------------
    wire    [1:0]   gtx8_rxpowerdown_i;
    wire    [1:0]   gtx8_txpowerdown_i;
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire    [1:0]   gtx8_rxchariscomma_i;
    wire    [1:0]   gtx8_rxcharisk_i;
    wire    [1:0]   gtx8_rxdisperr_i;
    wire    [1:0]   gtx8_rxnotintable_i;
    //----------------- Receive Ports - Clock Correction Ports -----------------
    wire    [2:0]   gtx8_rxclkcorcnt_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            gtx8_rxbyterealign_i;
    wire            gtx8_rxcommadet_i;
    wire            gtx8_rxenmcommaalign_i;
    wire            gtx8_rxenpcommaalign_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [15:0]  gtx8_rxdata_i;
    wire            gtx8_rxreset_i;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    wire            gtx8_rxcdrreset_i;
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    wire    [2:0]   gtx8_rxbufstatus_i;
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    wire    [1:0]   gtx8_rxlossofsync_i;
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    wire            gtx8_gtxrxreset_i;
    wire            gtx8_pllrxreset_i;
    wire            gtx8_rxplllkdet_i;
    wire            gtx8_rxresetdone_i;
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    wire            gtx8_rxvalid_i;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    wire            gtx8_rxpolarity_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [15:0]  gtx8_txdata_i;
    wire            gtx8_txoutclk_i;
    wire            gtx8_txreset_i;
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    wire            gtx8_txdlyaligndisable_i;
    wire            gtx8_txdlyalignmonenb_i;
    wire    [7:0]   gtx8_txdlyalignmonitor_i;
    wire            gtx8_txdlyalignreset_i;
    wire            gtx8_txenpmaphasealign_i;
    wire            gtx8_txpmasetphase_i;
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    wire            gtx8_gtxtxreset_i;
    wire            gtx8_txresetdone_i;


    //________________________________________________________________________
    //________________________________________________________________________
    //GTX9   (X0Y9)

    //---------------------- Loopback and Powerdown Ports ----------------------
    wire    [1:0]   gtx9_rxpowerdown_i;
    wire    [1:0]   gtx9_txpowerdown_i;
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire    [1:0]   gtx9_rxchariscomma_i;
    wire    [1:0]   gtx9_rxcharisk_i;
    wire    [1:0]   gtx9_rxdisperr_i;
    wire    [1:0]   gtx9_rxnotintable_i;
    //----------------- Receive Ports - Clock Correction Ports -----------------
    wire    [2:0]   gtx9_rxclkcorcnt_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            gtx9_rxbyterealign_i;
    wire            gtx9_rxcommadet_i;
    wire            gtx9_rxenmcommaalign_i;
    wire            gtx9_rxenpcommaalign_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [15:0]  gtx9_rxdata_i;
    wire            gtx9_rxreset_i;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    wire            gtx9_rxcdrreset_i;
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    wire    [2:0]   gtx9_rxbufstatus_i;
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    wire    [1:0]   gtx9_rxlossofsync_i;
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    wire            gtx9_gtxrxreset_i;
    wire            gtx9_pllrxreset_i;
    wire            gtx9_rxplllkdet_i;
    wire            gtx9_rxresetdone_i;
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    wire            gtx9_rxvalid_i;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    wire            gtx9_rxpolarity_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [15:0]  gtx9_txdata_i;
    wire            gtx9_txoutclk_i;
    wire            gtx9_txreset_i;
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    wire            gtx9_txdlyaligndisable_i;
    wire            gtx9_txdlyalignmonenb_i;
    wire    [7:0]   gtx9_txdlyalignmonitor_i;
    wire            gtx9_txdlyalignreset_i;
    wire            gtx9_txenpmaphasealign_i;
    wire            gtx9_txpmasetphase_i;
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    wire            gtx9_gtxtxreset_i;
    wire            gtx9_txresetdone_i;


    //________________________________________________________________________
    //________________________________________________________________________
    //GTX10   (X0Y10)

    //---------------------- Loopback and Powerdown Ports ----------------------
    wire    [1:0]   gtx10_rxpowerdown_i;
    wire    [1:0]   gtx10_txpowerdown_i;
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire    [1:0]   gtx10_rxchariscomma_i;
    wire    [1:0]   gtx10_rxcharisk_i;
    wire    [1:0]   gtx10_rxdisperr_i;
    wire    [1:0]   gtx10_rxnotintable_i;
    //----------------- Receive Ports - Clock Correction Ports -----------------
    wire    [2:0]   gtx10_rxclkcorcnt_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            gtx10_rxbyterealign_i;
    wire            gtx10_rxcommadet_i;
    wire            gtx10_rxenmcommaalign_i;
    wire            gtx10_rxenpcommaalign_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [15:0]  gtx10_rxdata_i;
    wire            gtx10_rxreset_i;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    wire            gtx10_rxcdrreset_i;
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    wire    [2:0]   gtx10_rxbufstatus_i;
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    wire    [1:0]   gtx10_rxlossofsync_i;
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    wire            gtx10_gtxrxreset_i;
    wire            gtx10_pllrxreset_i;
    wire            gtx10_rxplllkdet_i;
    wire            gtx10_rxresetdone_i;
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    wire            gtx10_rxvalid_i;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    wire            gtx10_rxpolarity_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [15:0]  gtx10_txdata_i;
    wire            gtx10_txoutclk_i;
    wire            gtx10_txreset_i;
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    wire            gtx10_txdlyaligndisable_i;
    wire            gtx10_txdlyalignmonenb_i;
    wire    [7:0]   gtx10_txdlyalignmonitor_i;
    wire            gtx10_txdlyalignreset_i;
    wire            gtx10_txenpmaphasealign_i;
    wire            gtx10_txpmasetphase_i;
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    wire            gtx10_gtxtxreset_i;
    wire            gtx10_txresetdone_i;


    //________________________________________________________________________
    //________________________________________________________________________
    //GTX11   (X0Y11)

    //---------------------- Loopback and Powerdown Ports ----------------------
    wire    [1:0]   gtx11_rxpowerdown_i;
    wire    [1:0]   gtx11_txpowerdown_i;
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
    wire    [1:0]   gtx11_rxchariscomma_i;
    wire    [1:0]   gtx11_rxcharisk_i;
    wire    [1:0]   gtx11_rxdisperr_i;
    wire    [1:0]   gtx11_rxnotintable_i;
    //----------------- Receive Ports - Clock Correction Ports -----------------
    wire    [2:0]   gtx11_rxclkcorcnt_i;
    //------------- Receive Ports - Comma Detection and Alignment --------------
    wire            gtx11_rxbyterealign_i;
    wire            gtx11_rxcommadet_i;
    wire            gtx11_rxenmcommaalign_i;
    wire            gtx11_rxenpcommaalign_i;
    //----------------- Receive Ports - RX Data Path interface -----------------
    wire    [15:0]  gtx11_rxdata_i;
    wire            gtx11_rxreset_i;
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    wire            gtx11_rxcdrreset_i;
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
    wire    [2:0]   gtx11_rxbufstatus_i;
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    wire    [1:0]   gtx11_rxlossofsync_i;
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    wire            gtx11_gtxrxreset_i;
    wire            gtx11_pllrxreset_i;
    wire            gtx11_rxplllkdet_i;
    wire            gtx11_rxresetdone_i;
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    wire            gtx11_rxvalid_i;
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    wire            gtx11_rxpolarity_i;
    //---------------- Transmit Ports - TX Data Path interface -----------------
    wire    [15:0]  gtx11_txdata_i;
    wire            gtx11_txoutclk_i;
    wire            gtx11_txreset_i;
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    wire            gtx11_txdlyaligndisable_i;
    wire            gtx11_txdlyalignmonenb_i;
    wire    [7:0]   gtx11_txdlyalignmonitor_i;
    wire            gtx11_txdlyalignreset_i;
    wire            gtx11_txenpmaphasealign_i;
    wire            gtx11_txpmasetphase_i;
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    wire            gtx11_gtxtxreset_i;
    wire            gtx11_txresetdone_i;




    //----------------------------- Global Signals -----------------------------
    wire            gtx0_tx_system_reset_c;
    wire            gtx0_rx_system_reset_c;
    wire            gtx1_tx_system_reset_c;
    wire            gtx1_rx_system_reset_c;
    wire            gtx2_tx_system_reset_c;
    wire            gtx2_rx_system_reset_c;
    wire            gtx3_tx_system_reset_c;
    wire            gtx3_rx_system_reset_c;
    wire            gtx4_tx_system_reset_c;
    wire            gtx4_rx_system_reset_c;
    wire            gtx5_tx_system_reset_c;
    wire            gtx5_rx_system_reset_c;
    wire            gtx6_tx_system_reset_c;
    wire            gtx6_rx_system_reset_c;
    wire            gtx7_tx_system_reset_c;
    wire            gtx7_rx_system_reset_c;
    wire            gtx8_tx_system_reset_c;
    wire            gtx8_rx_system_reset_c;
    wire            gtx9_tx_system_reset_c;
    wire            gtx9_rx_system_reset_c;
    wire            gtx10_tx_system_reset_c;
    wire            gtx10_rx_system_reset_c;
    wire            gtx11_tx_system_reset_c;
    wire            gtx11_rx_system_reset_c;
    wire            tied_to_ground_i;
    wire    [63:0]  tied_to_ground_vec_i;
    wire            tied_to_vcc_i;
    wire    [7:0]   tied_to_vcc_vec_i;
    wire            drp_clk_in_i;

    //--------------------------- User Clocks ---------------------------------
//    wire            snap_clk2;


    //--------------------------- Reference Clocks ----------------------------
    
    wire            q1_clk1_refclk_i;
    wire            q1_clk1_refclk_i_bufg;
    //--------------------- Frame check/gen Module Signals --------------------
    wire            gtx0_matchn_i;
    
    wire    [23:0]  gtx0_txdata_float_i;
    
    
    wire            gtx0_block_sync_i;
    wire            gtx0_track_data_i;
    wire    [7:0]   gtx0_error_count_i;
    wire            gtx0_frame_check_reset_i;
    wire            gtx0_inc_in_i;
    wire            gtx0_inc_out_i;
    wire    [15:0]  gtx0_unscrambled_data_i;

    wire            gtx1_matchn_i;
    
    wire    [23:0]  gtx1_txdata_float_i;
    
    
    wire            gtx1_block_sync_i;
    wire            gtx1_track_data_i;
    wire    [7:0]   gtx1_error_count_i;
    wire            gtx1_frame_check_reset_i;
    wire            gtx1_inc_in_i;
    wire            gtx1_inc_out_i;
    wire    [15:0]  gtx1_unscrambled_data_i;

    wire            gtx2_matchn_i;
    
    wire    [23:0]  gtx2_txdata_float_i;
    
    
    wire            gtx2_block_sync_i;
    wire            gtx2_track_data_i;
    wire    [7:0]   gtx2_error_count_i;
    wire            gtx2_frame_check_reset_i;
    wire            gtx2_inc_in_i;
    wire            gtx2_inc_out_i;
    wire    [15:0]  gtx2_unscrambled_data_i;

    wire            gtx3_matchn_i;
    
    wire    [23:0]  gtx3_txdata_float_i;
    
    
    wire            gtx3_block_sync_i;
    wire            gtx3_track_data_i;
    wire    [7:0]   gtx3_error_count_i;
    wire            gtx3_frame_check_reset_i;
    wire            gtx3_inc_in_i;
    wire            gtx3_inc_out_i;
    wire    [15:0]  gtx3_unscrambled_data_i;

    wire            gtx4_matchn_i;
    
    wire    [23:0]  gtx4_txdata_float_i;
    
    
    wire            gtx4_block_sync_i;
    wire            gtx4_track_data_i;
    wire    [7:0]   gtx4_error_count_i;
    wire            gtx4_frame_check_reset_i;
    wire            gtx4_inc_in_i;
    wire            gtx4_inc_out_i;
    wire    [15:0]  gtx4_unscrambled_data_i;

    wire            gtx5_matchn_i;
    
    wire    [23:0]  gtx5_txdata_float_i;
    
    
    wire            gtx5_block_sync_i;
    wire            gtx5_track_data_i;
    wire    [7:0]   gtx5_error_count_i;
    wire            gtx5_frame_check_reset_i;
    wire            gtx5_inc_in_i;
    wire            gtx5_inc_out_i;
    wire    [15:0]  gtx5_unscrambled_data_i;

    wire            gtx6_matchn_i;
    
    wire    [23:0]  gtx6_txdata_float_i;
    
    
    wire            gtx6_block_sync_i;
    wire            gtx6_track_data_i;
    wire    [7:0]   gtx6_error_count_i;
    wire            gtx6_frame_check_reset_i;
    wire            gtx6_inc_in_i;
    wire            gtx6_inc_out_i;
    wire    [15:0]  gtx6_unscrambled_data_i;

    wire            gtx7_matchn_i;
    
    wire    [23:0]  gtx7_txdata_float_i;
    
    
    wire            gtx7_block_sync_i;
    wire            gtx7_track_data_i;
    wire    [7:0]   gtx7_error_count_i;
    wire            gtx7_frame_check_reset_i;
    wire            gtx7_inc_in_i;
    wire            gtx7_inc_out_i;
    wire    [15:0]  gtx7_unscrambled_data_i;

    wire            gtx8_matchn_i;
    
    wire    [23:0]  gtx8_txdata_float_i;
    
    
    wire            gtx8_block_sync_i;
    wire            gtx8_track_data_i;
    wire    [7:0]   gtx8_error_count_i;
    wire            gtx8_frame_check_reset_i;
    wire            gtx8_inc_in_i;
    wire            gtx8_inc_out_i;
    wire    [15:0]  gtx8_unscrambled_data_i;

    wire            gtx9_matchn_i;
    
    wire    [23:0]  gtx9_txdata_float_i;
    
    
    wire            gtx9_block_sync_i;
    wire            gtx9_track_data_i;
    wire    [7:0]   gtx9_error_count_i;
    wire            gtx9_frame_check_reset_i;
    wire            gtx9_inc_in_i;
    wire            gtx9_inc_out_i;
    wire    [15:0]  gtx9_unscrambled_data_i;

    wire            gtx10_matchn_i;
    
    wire    [23:0]  gtx10_txdata_float_i;
    
    
    wire            gtx10_block_sync_i;
    wire            gtx10_track_data_i;
    wire    [7:0]   gtx10_error_count_i;
    wire            gtx10_frame_check_reset_i;
    wire            gtx10_inc_in_i;
    wire            gtx10_inc_out_i;
    wire    [15:0]  gtx10_unscrambled_data_i;

    wire            gtx11_matchn_i;
    
    wire    [23:0]  gtx11_txdata_float_i;
    
    
    wire            gtx11_block_sync_i;
    wire            gtx11_track_data_i;
    wire    [7:0]   gtx11_error_count_i;
    wire            gtx11_frame_check_reset_i;
    wire            gtx11_inc_in_i;
    wire            gtx11_inc_out_i;
    wire    [15:0]  gtx11_unscrambled_data_i;

    wire            reset_on_data_error_i;
    wire            track_data_out_i;

    //----------------------- Sync Module Signals -----------------------------


    wire            gtx0_tx_sync_done_i;
    wire            gtx0_reset_txsync_c;
    wire            gtx1_tx_sync_done_i;
    wire            gtx1_reset_txsync_c;
    wire            gtx2_tx_sync_done_i;
    wire            gtx2_reset_txsync_c;
    wire            gtx3_tx_sync_done_i;
    wire            gtx3_reset_txsync_c;
    wire            gtx4_tx_sync_done_i;
    wire            gtx4_reset_txsync_c;
    wire            gtx5_tx_sync_done_i;
    wire            gtx5_reset_txsync_c;
    wire            gtx6_tx_sync_done_i;
    wire            gtx6_reset_txsync_c;
    wire            gtx7_tx_sync_done_i;
    wire            gtx7_reset_txsync_c;
    wire            gtx8_tx_sync_done_i;
    wire            gtx8_reset_txsync_c;
    wire            gtx9_tx_sync_done_i;
    wire            gtx9_reset_txsync_c;
    wire            gtx10_tx_sync_done_i;
    wire            gtx10_reset_txsync_c;
    wire            gtx11_tx_sync_done_i;
    wire            gtx11_reset_txsync_c;

    wire            gtxtxreset_i;
    wire            gtxrxreset_i;
    wire    [3:0]   mux_sel_i;

    wire            user_tx_reset_i;
    wire            user_rx_reset_i;

//**************************** Main Body of Code *******************************

    //  Static signal Assigments    
    assign tied_to_ground_i             = 1'b0;
    assign tied_to_ground_vec_i         = 64'h0000000000000000;
    assign tied_to_vcc_i                = 1'b1;
    assign tied_to_vcc_vec_i            = 8'hff;

    assign rxdv_diff[0] = rxdv_snapr[0]^gtx0_rxvalid_i;
    assign rxdv_diff[1] = rxdv_snapr[1]^gtx1_rxvalid_i;
    assign rxdv_diff[2] = rxdv_snapr[2]^gtx2_rxvalid_i;
    assign rxdv_diff[3] = rxdv_snapr[3]^gtx3_rxvalid_i;
    assign rxdv_diff[4] = rxdv_snapr[4]^gtx8_rxvalid_i;
    assign rxdv_diff[5] = rxdv_snapr[5]^gtx9_rxvalid_i;
    assign rxdv_diff[6] = rxdv_snapr[6]^gtx10_rxvalid_i;
    assign rxdv_diff[7] = rxdv_snapr[7]^gtx11_rxvalid_i;
    assign rxcomma_diff[0] = rxcomma_snapr[0]^gtx0_rxcommadet_i;
    assign rxcomma_diff[1] = rxcomma_snapr[1]^gtx1_rxcommadet_i;
    assign rxcomma_diff[2] = rxcomma_snapr[2]^gtx2_rxcommadet_i;
    assign rxcomma_diff[3] = rxcomma_snapr[3]^gtx3_rxcommadet_i;
    assign rxcomma_diff[4] = rxcomma_snapr[4]^gtx8_rxcommadet_i;
    assign rxcomma_diff[5] = rxcomma_snapr[5]^gtx9_rxcommadet_i;
    assign rxcomma_diff[6] = rxcomma_snapr[6]^gtx10_rxcommadet_i;
    assign rxcomma_diff[7] = rxcomma_snapr[7]^gtx11_rxcommadet_i;



    //---------------------Dedicated GTX Reference Clock Inputs ---------------
    // The dedicated reference clock inputs you selected in the GUI are implemented using
    // IBUFDS_GTXE1 instances.
    //
    // In the UCF file for this example design, you will see that each of
    // these IBUFDS_GTXE1 instances has been LOCed to a particular set of pins. By LOCing to these
    // locations, we tell the tools to use the dedicated input buffers to the GTX reference
    // clock network, rather than general purpose IOs. To select other pins, consult the 
    // Implementation chapter of UG___, or rerun the wizard.
    //
    // This network is the highest performace (lowest jitter) option for providing clocks
    // to the GTX transceivers.
    
    IBUFDS_GTXE1 q1_clk1_refclk_ibufds_i
    (
        .O                              (q1_clk1_refclk_i),
        .ODIV2                          (),
        .CEB                            (tied_to_ground_i),
        .I                              (ck_160p),
        .IB                             (ck_160n)
    );

 
    

    BUFG q1_clk1_refclk_bufg_i
    (
        .I                              (q1_clk1_refclk_i),
        .O                              (q1_clk1_refclk_i_bufg)
    );



    //--------------------------------- User Clocks ---------------------------
    
    // The clock resources in this section were added based on userclk source selections on
    // the Latency, Buffering, and Clocking page of the GUI. A few notes about user clocks:
    // * The userclk and userclk2 for each GTX datapath (TX and RX) must be phase aligned to 
    //   avoid data errors in the fabric interface whenever the datapath is wider than 10 bits
    // * To minimize clock resources, you can share clocks between GTXs. GTXs using the same frequency
    //   or multiples of the same frequency can be accomadated using MMCMs. Use caution when
    //   using RXRECCLK as a clock source, however - these clocks can typically only be shared if all
    //   the channels using the clock are receiving data from TX channels that share a reference clock 
    //   source with each other.

    BUFG txoutclk_bufg0_i
    (
        .I                              (gtx3_txoutclk_i),
        .O                              (snap_clk2)
    );

   assign ck_160_plllkdet = gtx3_rxplllkdet_i;






    //--------------------------- The GTX Wrapper -----------------------------
    
    // Use the instantiation template in the example directory to add the GTX wrapper to your design.
    // In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    // checker. The GTXs will reset, then attempt to align and transmit data. If channel bonding is 
    // enabled, bonding should occur after alignment.
    
    SNAP12_T20R20 #
    (
        .WRAPPER_SIM_GTXRESET_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP)
    )
    snap12_t20r20_i
    (
        //_____________________________________________________________________
        //_____________________________________________________________________
        .gtx_wait   (gtx_wait),
        .rxdv_snapr (rxdv_snapr),
        .rxcomma_snapr   (rxcomma_snapr),
        .check_ok_snapr  (check_ok_snapr),
        .check_bad_snapr (check_bad_snapr),
        .good_byte (good_byte),
        .bad_byte  (bad_byte),
        .lost_byte (lost_byte),
        .errcount0 (snap_err0),
        .errcount1 (snap_err1),
        .errcount2 (snap_err2),
        .errcount3 (snap_err3),
        .errcount4 (snap_err4),
        .errcount5 (snap_err5),
        .errcount6 (snap_err6),
        .errcount7 (snap_err7),
        .GTXi_RXDATA_OUT (rxdata_i),  // the one select gtx data to monitor...
        .GTXi_RXK_OUT (RXK_OUT),      // the K that goes with it
//
        //GTX0  (X0Y0)
        //---------------------- Loopback and Powerdown Ports ----------------------
//jg        .GTX0_RXPOWERDOWN_IN            (gtx0_rxpowerdown_i),
//jg        .GTX0_TXPOWERDOWN_IN            (gtx0_txpowerdown_i),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .GTX0_RXCLKCORCNT_OUT           (gtx0_rxclkcorcnt_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .GTX0_RXBYTEREALIGN_OUT         (gtx0_rxbyterealign_i),
        .GTX0_RXCOMMADET_OUT            (gtx0_rxcommadet_i),    //jg: useful?
        .GTX0_RXENMCOMMAALIGN_IN        (snap_commaalign),
        .GTX0_RXENPCOMMAALIGN_IN        (snap_commaalign),
        //----------------- Receive Ports - RX Data Path interface -----------------
//jg        .GTX0_RXDATA_OUT                (gtx0_rxdata_i),
        .GTX0_RXRESET_IN                (!ck_160_plllkdet),
        .GTX0_RXUSRCLK2_IN              (snap_clk2),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .GTX0_RXCDRRESET_IN             (gtx0_rxcdrreset_i),
        .GTX0_RXN_IN                    (RXN[0]),
        .GTX0_RXP_IN                    (RXP[0]),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .GTX0_RXLOSSOFSYNC_OUT          (gtx0_rxlossofsync_i),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTX0_GTXRXRESET_IN             (gtx0_gtxrxreset_i),
        .GTX0_MGTREFCLKRX_IN            (q1_clk1_refclk_i),
        .GTX0_PLLRXRESET_IN             (gtx0_pllrxreset_i),
        .GTX0_RXPLLLKDET_OUT            (gtx0_rxplllkdet_i),
        .GTX0_RXRESETDONE_OUT           (gtx0_rxresetdone_i),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .GTX0_RXVALID_OUT               (gtx0_rxvalid_i),       //jg: useful?
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .GTX0_RXPOLARITY_IN             (gtx0_rxpolarity_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GTX0_SEED_IN                 (),
        .GTX0_RXSEED                  (seed_in[0]),
        .GTX0_TXOUTCLK_OUT              (gtx0_txoutclk_i),
        .GTX0_TXRESET_IN                (!ck_160_plllkdet),
        .GTX0_TXUSRCLK2_IN              (snap_clk2),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GTX0_TXN_OUT                   (),
        .GTX0_TXP_OUT                   (),
        .gtx0_force_error               (),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .GTX0_TXDLYALIGNDISABLE_IN      (gtx0_txdlyaligndisable_i),
        .GTX0_TXDLYALIGNMONENB_IN       (gtx0_txdlyalignmonenb_i),
        .GTX0_TXDLYALIGNMONITOR_OUT     (gtx0_txdlyalignmonitor_i),
        .GTX0_TXDLYALIGNRESET_IN        (gtx0_txdlyalignreset_i),
        .GTX0_TXENPMAPHASEALIGN_IN      (gtx0_txenpmaphasealign_i),
        .GTX0_TXPMASETPHASE_IN          (gtx0_txpmasetphase_i),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTX0_GTXTXRESET_IN             (gtx0_gtxtxreset_i),
        .GTX0_TXRESETDONE_OUT           (gtx0_txresetdone_i),


 
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GTX1  (X0Y1)
        //---------------------- Loopback and Powerdown Ports ----------------------
//jg        .GTX1_RXPOWERDOWN_IN            (gtx1_rxpowerdown_i),
//jg        .GTX1_TXPOWERDOWN_IN            (gtx1_txpowerdown_i),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .GTX1_RXCLKCORCNT_OUT           (gtx1_rxclkcorcnt_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .GTX1_RXBYTEREALIGN_OUT         (gtx1_rxbyterealign_i),
        .GTX1_RXCOMMADET_OUT            (gtx1_rxcommadet_i),
        .GTX1_RXENMCOMMAALIGN_IN        (snap_commaalign),
        .GTX1_RXENPCOMMAALIGN_IN        (snap_commaalign),
        //----------------- Receive Ports - RX Data Path interface -----------------
//jg        .GTX1_RXDATA_OUT                (gtx1_rxdata_i),
        .GTX1_RXRESET_IN                (!ck_160_plllkdet),
        .GTX1_RXUSRCLK2_IN              (snap_clk2),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .GTX1_RXCDRRESET_IN             (gtx1_rxcdrreset_i),
        .GTX1_RXN_IN                    (RXN[1]),
        .GTX1_RXP_IN                    (RXP[1]),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .GTX1_RXLOSSOFSYNC_OUT          (gtx1_rxlossofsync_i),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTX1_GTXRXRESET_IN             (gtx1_gtxrxreset_i),
        .GTX1_MGTREFCLKRX_IN            (q1_clk1_refclk_i),
        .GTX1_PLLRXRESET_IN             (gtx1_pllrxreset_i),
        .GTX1_RXPLLLKDET_OUT            (gtx1_rxplllkdet_i),
        .GTX1_RXRESETDONE_OUT           (gtx1_rxresetdone_i),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .GTX1_RXVALID_OUT               (gtx1_rxvalid_i),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .GTX1_RXPOLARITY_IN             (gtx1_rxpolarity_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GTX1_SEED_IN                 (),
        .GTX1_RXSEED                  (seed_in[1]),
        .GTX1_TXOUTCLK_OUT              (gtx1_txoutclk_i),
        .GTX1_TXRESET_IN                (!ck_160_plllkdet),
        .GTX1_TXUSRCLK2_IN              (snap_clk2),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GTX1_TXN_OUT                   (),
        .GTX1_TXP_OUT                   (),
        .gtx1_force_error               (),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .GTX1_TXDLYALIGNDISABLE_IN      (gtx1_txdlyaligndisable_i),
        .GTX1_TXDLYALIGNMONENB_IN       (gtx1_txdlyalignmonenb_i),
        .GTX1_TXDLYALIGNMONITOR_OUT     (gtx1_txdlyalignmonitor_i),
        .GTX1_TXDLYALIGNRESET_IN        (gtx1_txdlyalignreset_i),
        .GTX1_TXENPMAPHASEALIGN_IN      (gtx1_txenpmaphasealign_i),
        .GTX1_TXPMASETPHASE_IN          (gtx1_txpmasetphase_i),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTX1_GTXTXRESET_IN             (gtx1_gtxtxreset_i),
        .GTX1_TXRESETDONE_OUT           (gtx1_txresetdone_i),


 
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GTX2  (X0Y2)
        //---------------------- Loopback and Powerdown Ports ----------------------
//jg        .GTX2_RXPOWERDOWN_IN            (gtx2_rxpowerdown_i),
//jg        .GTX2_TXPOWERDOWN_IN            (gtx2_txpowerdown_i),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .GTX2_RXCLKCORCNT_OUT           (gtx2_rxclkcorcnt_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .GTX2_RXBYTEREALIGN_OUT         (gtx2_rxbyterealign_i),
        .GTX2_RXCOMMADET_OUT            (gtx2_rxcommadet_i),
        .GTX2_RXENMCOMMAALIGN_IN        (snap_commaalign),
        .GTX2_RXENPCOMMAALIGN_IN        (snap_commaalign),
        //----------------- Receive Ports - RX Data Path interface -----------------
//jg        .GTX2_RXDATA_OUT                (gtx2_rxdata_i),
        .GTX2_RXRESET_IN                (!ck_160_plllkdet),
        .GTX2_RXUSRCLK2_IN              (snap_clk2),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .GTX2_RXCDRRESET_IN             (gtx2_rxcdrreset_i),
        .GTX2_RXN_IN                    (RXN[2]),
        .GTX2_RXP_IN                    (RXP[2]),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .GTX2_RXLOSSOFSYNC_OUT          (gtx2_rxlossofsync_i),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTX2_GTXRXRESET_IN             (gtx2_gtxrxreset_i),
        .GTX2_MGTREFCLKRX_IN            (q1_clk1_refclk_i),
        .GTX2_PLLRXRESET_IN             (gtx2_pllrxreset_i),
        .GTX2_RXPLLLKDET_OUT            (gtx2_rxplllkdet_i),
        .GTX2_RXRESETDONE_OUT           (gtx2_rxresetdone_i),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .GTX2_RXVALID_OUT               (gtx2_rxvalid_i),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .GTX2_RXPOLARITY_IN             (gtx2_rxpolarity_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GTX2_SEED_IN                 (seed_in[7]),
        .GTX2_RXSEED                  (seed_in[2]),
        .GTX2_TXOUTCLK_OUT              (gtx2_txoutclk_i),
        .GTX2_TXRESET_IN                (!ck_160_plllkdet),
        .GTX2_TXUSRCLK2_IN              (snap_clk2),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GTX2_TXN_OUT                   (TXN[7]),
        .GTX2_TXP_OUT                   (TXP[7]),
        .gtx2_force_error               (force_err_wait & force_err_flag[7]),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .GTX2_TXDLYALIGNDISABLE_IN      (gtx2_txdlyaligndisable_i),
        .GTX2_TXDLYALIGNMONENB_IN       (gtx2_txdlyalignmonenb_i),
        .GTX2_TXDLYALIGNMONITOR_OUT     (gtx2_txdlyalignmonitor_i),
        .GTX2_TXDLYALIGNRESET_IN        (gtx2_txdlyalignreset_i),
        .GTX2_TXENPMAPHASEALIGN_IN      (gtx2_txenpmaphasealign_i),
        .GTX2_TXPMASETPHASE_IN          (gtx2_txpmasetphase_i),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTX2_GTXTXRESET_IN             (gtx2_gtxtxreset_i),
        .GTX2_TXRESETDONE_OUT           (gtx2_txresetdone_i),


 
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GTX3  (X0Y3)
        //---------------------- Loopback and Powerdown Ports ----------------------
//jg        .GTX3_RXPOWERDOWN_IN            (gtx3_rxpowerdown_i),
//jg        .GTX3_TXPOWERDOWN_IN            (gtx3_txpowerdown_i),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .GTX3_RXCLKCORCNT_OUT           (gtx3_rxclkcorcnt_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .GTX3_RXBYTEREALIGN_OUT         (gtx3_rxbyterealign_i),
        .GTX3_RXCOMMADET_OUT            (gtx3_rxcommadet_i),
        .GTX3_RXENMCOMMAALIGN_IN        (snap_commaalign),
        .GTX3_RXENPCOMMAALIGN_IN        (snap_commaalign),
        //----------------- Receive Ports - RX Data Path interface -----------------
//jg        .GTX3_RXDATA_OUT                (gtx3_rxdata_i),
        .GTX3_RXRESET_IN                (!ck_160_plllkdet),
        .GTX3_RXUSRCLK2_IN              (snap_clk2),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .GTX3_RXCDRRESET_IN             (gtx3_rxcdrreset_i),
        .GTX3_RXN_IN                    (RXN[3]),
        .GTX3_RXP_IN                    (RXP[3]),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .GTX3_RXLOSSOFSYNC_OUT          (gtx3_rxlossofsync_i),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTX3_GTXRXRESET_IN             (gtx3_gtxrxreset_i),
        .GTX3_MGTREFCLKRX_IN            (q1_clk1_refclk_i),
        .GTX3_PLLRXRESET_IN             (gtx3_pllrxreset_i),
        .GTX3_RXPLLLKDET_OUT            (gtx3_rxplllkdet_i),
        .GTX3_RXRESETDONE_OUT           (gtx3_rxresetdone_i),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .GTX3_RXVALID_OUT               (gtx3_rxvalid_i),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .GTX3_RXPOLARITY_IN             (gtx3_rxpolarity_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GTX3_SEED_IN                 (seed_in[0]),
        .GTX3_RXSEED                  (seed_in[3]),
        .GTX3_TXOUTCLK_OUT              (gtx3_txoutclk_i),
        .GTX3_TXRESET_IN                (!ck_160_plllkdet),
        .GTX3_TXUSRCLK2_IN              (snap_clk2),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GTX3_TXN_OUT                   (TXN[0]),
        .GTX3_TXP_OUT                   (TXP[0]),
        .gtx3_force_error               (force_err_wait & force_err_flag[0]),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .GTX3_TXDLYALIGNDISABLE_IN      (gtx3_txdlyaligndisable_i),
        .GTX3_TXDLYALIGNMONENB_IN       (gtx3_txdlyalignmonenb_i),
        .GTX3_TXDLYALIGNMONITOR_OUT     (gtx3_txdlyalignmonitor_i),
        .GTX3_TXDLYALIGNRESET_IN        (gtx3_txdlyalignreset_i),
        .GTX3_TXENPMAPHASEALIGN_IN      (gtx3_txenpmaphasealign_i),
        .GTX3_TXPMASETPHASE_IN          (gtx3_txpmasetphase_i),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTX3_GTXTXRESET_IN             (gtx3_gtxtxreset_i),
        .GTX3_TXRESETDONE_OUT           (gtx3_txresetdone_i),


 
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GTX4  (X0Y4)
        //---------------------- Loopback and Powerdown Ports ----------------------
//jg        .GTX4_RXPOWERDOWN_IN            (gtx4_rxpowerdown_i),
//jg        .GTX4_TXPOWERDOWN_IN            (gtx4_txpowerdown_i),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .GTX4_RXCLKCORCNT_OUT           (gtx4_rxclkcorcnt_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .GTX4_RXBYTEREALIGN_OUT         (gtx4_rxbyterealign_i),
        .GTX4_RXCOMMADET_OUT            (gtx4_rxcommadet_i),
        .GTX4_RXENMCOMMAALIGN_IN        (snap_commaalign),
        .GTX4_RXENPCOMMAALIGN_IN        (snap_commaalign),
        //----------------- Receive Ports - RX Data Path interface -----------------
//jg        .GTX4_RXDATA_OUT                (gtx4_rxdata_i),
        .GTX4_RXRESET_IN                (!ck_160_plllkdet),
        .GTX4_RXUSRCLK2_IN              (snap_clk2),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .GTX4_RXCDRRESET_IN             (gtx4_rxcdrreset_i),
        .GTX4_RXN_IN                    (),
        .GTX4_RXP_IN                    (),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .GTX4_RXLOSSOFSYNC_OUT          (gtx4_rxlossofsync_i),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTX4_GTXRXRESET_IN             (gtx4_gtxrxreset_i),
        .GTX4_MGTREFCLKRX_IN            (q1_clk1_refclk_i),
        .GTX4_PLLRXRESET_IN             (gtx4_pllrxreset_i),
        .GTX4_RXPLLLKDET_OUT            (gtx4_rxplllkdet_i),
        .GTX4_RXRESETDONE_OUT           (gtx4_rxresetdone_i),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .GTX4_RXVALID_OUT               (gtx4_rxvalid_i),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .GTX4_RXPOLARITY_IN             (gtx4_rxpolarity_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GTX4_SEED_IN                 (seed_in[1]),
        .GTX4_RXSEED                  (seed_in[0]),
        .GTX4_TXOUTCLK_OUT              (gtx4_txoutclk_i),
        .GTX4_TXRESET_IN                (!ck_160_plllkdet),
        .GTX4_TXUSRCLK2_IN              (snap_clk2),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GTX4_TXN_OUT                   (TXN[1]),
        .GTX4_TXP_OUT                   (TXP[1]),
        .gtx4_force_error               (force_err_wait & force_err_flag[1]),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .GTX4_TXDLYALIGNDISABLE_IN      (gtx4_txdlyaligndisable_i),
        .GTX4_TXDLYALIGNMONENB_IN       (gtx4_txdlyalignmonenb_i),
        .GTX4_TXDLYALIGNMONITOR_OUT     (gtx4_txdlyalignmonitor_i),
        .GTX4_TXDLYALIGNRESET_IN        (gtx4_txdlyalignreset_i),
        .GTX4_TXENPMAPHASEALIGN_IN      (gtx4_txenpmaphasealign_i),
        .GTX4_TXPMASETPHASE_IN          (gtx4_txpmasetphase_i),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTX4_GTXTXRESET_IN             (gtx4_gtxtxreset_i),
        .GTX4_TXRESETDONE_OUT           (gtx4_txresetdone_i),


 
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GTX5  (X0Y5)
        //---------------------- Loopback and Powerdown Ports ----------------------
//jg        .GTX5_RXPOWERDOWN_IN            (gtx5_rxpowerdown_i),
//jg        .GTX5_TXPOWERDOWN_IN            (gtx5_txpowerdown_i),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .GTX5_RXCLKCORCNT_OUT           (gtx5_rxclkcorcnt_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .GTX5_RXBYTEREALIGN_OUT         (gtx5_rxbyterealign_i),
        .GTX5_RXCOMMADET_OUT            (gtx5_rxcommadet_i),
        .GTX5_RXENMCOMMAALIGN_IN        (snap_commaalign),
        .GTX5_RXENPCOMMAALIGN_IN        (snap_commaalign),
        //----------------- Receive Ports - RX Data Path interface -----------------
//jg        .GTX5_RXDATA_OUT                (gtx5_rxdata_i),
        .GTX5_RXRESET_IN                (!ck_160_plllkdet),
        .GTX5_RXUSRCLK2_IN              (snap_clk2),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .GTX5_RXCDRRESET_IN             (gtx5_rxcdrreset_i),
        .GTX5_RXN_IN                    (),
        .GTX5_RXP_IN                    (),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .GTX5_RXLOSSOFSYNC_OUT          (gtx5_rxlossofsync_i),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTX5_GTXRXRESET_IN             (gtx5_gtxrxreset_i),
        .GTX5_MGTREFCLKRX_IN            (q1_clk1_refclk_i),
        .GTX5_PLLRXRESET_IN             (gtx5_pllrxreset_i),
        .GTX5_RXPLLLKDET_OUT            (gtx5_rxplllkdet_i),
        .GTX5_RXRESETDONE_OUT           (gtx5_rxresetdone_i),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .GTX5_RXVALID_OUT               (gtx5_rxvalid_i),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .GTX5_RXPOLARITY_IN             (gtx5_rxpolarity_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GTX5_SEED_IN                 (),
        .GTX5_RXSEED                  (seed_in[1]),
        .GTX5_TXOUTCLK_OUT              (gtx5_txoutclk_i),
        .GTX5_TXRESET_IN                (!ck_160_plllkdet),
        .GTX5_TXUSRCLK2_IN              (snap_clk2),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GTX5_TXN_OUT                   (),
        .GTX5_TXP_OUT                   (),
        .gtx5_force_error               (),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .GTX5_TXDLYALIGNDISABLE_IN      (gtx5_txdlyaligndisable_i),
        .GTX5_TXDLYALIGNMONENB_IN       (gtx5_txdlyalignmonenb_i),
        .GTX5_TXDLYALIGNMONITOR_OUT     (gtx5_txdlyalignmonitor_i),
        .GTX5_TXDLYALIGNRESET_IN        (gtx5_txdlyalignreset_i),
        .GTX5_TXENPMAPHASEALIGN_IN      (gtx5_txenpmaphasealign_i),
        .GTX5_TXPMASETPHASE_IN          (gtx5_txpmasetphase_i),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTX5_GTXTXRESET_IN             (gtx5_gtxtxreset_i),
        .GTX5_TXRESETDONE_OUT           (gtx5_txresetdone_i),


 
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GTX6  (X0Y6)
        //---------------------- Loopback and Powerdown Ports ----------------------
//jg        .GTX6_RXPOWERDOWN_IN            (gtx6_rxpowerdown_i),
//jg        .GTX6_TXPOWERDOWN_IN            (gtx6_txpowerdown_i),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .GTX6_RXCLKCORCNT_OUT           (gtx6_rxclkcorcnt_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .GTX6_RXBYTEREALIGN_OUT         (gtx6_rxbyterealign_i),
        .GTX6_RXCOMMADET_OUT            (gtx6_rxcommadet_i),
        .GTX6_RXENMCOMMAALIGN_IN        (snap_commaalign),
        .GTX6_RXENPCOMMAALIGN_IN        (snap_commaalign),
        //----------------- Receive Ports - RX Data Path interface -----------------
//jg        .GTX6_RXDATA_OUT                (gtx6_rxdata_i),
        .GTX6_RXRESET_IN                (!ck_160_plllkdet),
        .GTX6_RXUSRCLK2_IN              (snap_clk2),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .GTX6_RXCDRRESET_IN             (gtx6_rxcdrreset_i),
        .GTX6_RXN_IN                    (),
        .GTX6_RXP_IN                    (),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .GTX6_RXLOSSOFSYNC_OUT          (gtx6_rxlossofsync_i),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTX6_GTXRXRESET_IN             (gtx6_gtxrxreset_i),
        .GTX6_MGTREFCLKRX_IN            (q1_clk1_refclk_i),
        .GTX6_PLLRXRESET_IN             (gtx6_pllrxreset_i),
        .GTX6_RXPLLLKDET_OUT            (gtx6_rxplllkdet_i),
        .GTX6_RXRESETDONE_OUT           (gtx6_rxresetdone_i),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .GTX6_RXVALID_OUT               (gtx6_rxvalid_i),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .GTX6_RXPOLARITY_IN             (gtx6_rxpolarity_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GTX6_SEED_IN                 (),
        .GTX6_RXSEED                  (seed_in[2]),
        .GTX6_TXOUTCLK_OUT              (gtx6_txoutclk_i),
        .GTX6_TXRESET_IN                (!ck_160_plllkdet),
        .GTX6_TXUSRCLK2_IN              (snap_clk2),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GTX6_TXN_OUT                   (),
        .GTX6_TXP_OUT                   (),
        .gtx6_force_error               (),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .GTX6_TXDLYALIGNDISABLE_IN      (gtx6_txdlyaligndisable_i),
        .GTX6_TXDLYALIGNMONENB_IN       (gtx6_txdlyalignmonenb_i),
        .GTX6_TXDLYALIGNMONITOR_OUT     (gtx6_txdlyalignmonitor_i),
        .GTX6_TXDLYALIGNRESET_IN        (gtx6_txdlyalignreset_i),
        .GTX6_TXENPMAPHASEALIGN_IN      (gtx6_txenpmaphasealign_i),
        .GTX6_TXPMASETPHASE_IN          (gtx6_txpmasetphase_i),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTX6_GTXTXRESET_IN             (gtx6_gtxtxreset_i),
        .GTX6_TXRESETDONE_OUT           (gtx6_txresetdone_i),


 
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GTX7  (X0Y7)
        //---------------------- Loopback and Powerdown Ports ----------------------
//jg        .GTX7_RXPOWERDOWN_IN            (gtx7_rxpowerdown_i),
//jg        .GTX7_TXPOWERDOWN_IN            (gtx7_txpowerdown_i),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .GTX7_RXCLKCORCNT_OUT           (gtx7_rxclkcorcnt_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .GTX7_RXBYTEREALIGN_OUT         (gtx7_rxbyterealign_i),
        .GTX7_RXCOMMADET_OUT            (gtx7_rxcommadet_i),
        .GTX7_RXENMCOMMAALIGN_IN        (snap_commaalign),
        .GTX7_RXENPCOMMAALIGN_IN        (snap_commaalign),
        //----------------- Receive Ports - RX Data Path interface -----------------
//jg        .GTX7_RXDATA_OUT                (gtx7_rxdata_i),
        .GTX7_RXRESET_IN                (!ck_160_plllkdet),
        .GTX7_RXUSRCLK2_IN              (snap_clk2),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .GTX7_RXCDRRESET_IN             (gtx7_rxcdrreset_i),
        .GTX7_RXN_IN                    (),
        .GTX7_RXP_IN                    (),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .GTX7_RXLOSSOFSYNC_OUT          (gtx7_rxlossofsync_i),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTX7_GTXRXRESET_IN             (gtx7_gtxrxreset_i),
        .GTX7_MGTREFCLKRX_IN            (q1_clk1_refclk_i),
        .GTX7_PLLRXRESET_IN             (gtx7_pllrxreset_i),
        .GTX7_RXPLLLKDET_OUT            (gtx7_rxplllkdet_i),
        .GTX7_RXRESETDONE_OUT           (gtx7_rxresetdone_i),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .GTX7_RXVALID_OUT               (gtx7_rxvalid_i),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .GTX7_RXPOLARITY_IN             (gtx7_rxpolarity_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GTX7_SEED_IN                 (seed_in[2]),
        .GTX7_RXSEED                  (seed_in[3]),
        .GTX7_TXOUTCLK_OUT              (gtx7_txoutclk_i),
        .GTX7_TXRESET_IN                (!ck_160_plllkdet),
        .GTX7_TXUSRCLK2_IN              (snap_clk2),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GTX7_TXN_OUT                   (TXN[2]),
        .GTX7_TXP_OUT                   (TXP[2]),
        .gtx7_force_error               (force_err_wait & force_err_flag[2]),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .GTX7_TXDLYALIGNDISABLE_IN      (gtx7_txdlyaligndisable_i),
        .GTX7_TXDLYALIGNMONENB_IN       (gtx7_txdlyalignmonenb_i),
        .GTX7_TXDLYALIGNMONITOR_OUT     (gtx7_txdlyalignmonitor_i),
        .GTX7_TXDLYALIGNRESET_IN        (gtx7_txdlyalignreset_i),
        .GTX7_TXENPMAPHASEALIGN_IN      (gtx7_txenpmaphasealign_i),
        .GTX7_TXPMASETPHASE_IN          (gtx7_txpmasetphase_i),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTX7_GTXTXRESET_IN             (gtx7_gtxtxreset_i),
        .GTX7_TXRESETDONE_OUT           (gtx7_txresetdone_i),


 
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GTX8  (X0Y8)
        //---------------------- Loopback and Powerdown Ports ----------------------
//jg        .GTX8_RXPOWERDOWN_IN            (gtx8_rxpowerdown_i),
//jg        .GTX8_TXPOWERDOWN_IN            (gtx8_txpowerdown_i),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .GTX8_RXCLKCORCNT_OUT           (gtx8_rxclkcorcnt_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .GTX8_RXBYTEREALIGN_OUT         (gtx8_rxbyterealign_i),
        .GTX8_RXCOMMADET_OUT            (gtx8_rxcommadet_i),
        .GTX8_RXENMCOMMAALIGN_IN        (snap_commaalign),
        .GTX8_RXENPCOMMAALIGN_IN        (snap_commaalign),
        //----------------- Receive Ports - RX Data Path interface -----------------
//jg        .GTX8_RXDATA_OUT                (gtx8_rxdata_i),
        .GTX8_RXRESET_IN                (!ck_160_plllkdet),
        .GTX8_RXUSRCLK2_IN              (snap_clk2),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .GTX8_RXCDRRESET_IN             (gtx8_rxcdrreset_i),
        .GTX8_RXN_IN                    (RXN[4]),
        .GTX8_RXP_IN                    (RXP[4]),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .GTX8_RXLOSSOFSYNC_OUT          (gtx8_rxlossofsync_i),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTX8_GTXRXRESET_IN             (gtx8_gtxrxreset_i),
        .GTX8_MGTREFCLKRX_IN            (q1_clk1_refclk_i),
        .GTX8_PLLRXRESET_IN             (gtx8_pllrxreset_i),
        .GTX8_RXPLLLKDET_OUT            (gtx8_rxplllkdet_i),
        .GTX8_RXRESETDONE_OUT           (gtx8_rxresetdone_i),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .GTX8_RXVALID_OUT               (gtx8_rxvalid_i),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .GTX8_RXPOLARITY_IN             (gtx8_rxpolarity_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GTX8_SEED_IN                 (seed_in[3]),
        .GTX8_RXSEED                  (seed_in[4]),
        .GTX8_TXOUTCLK_OUT              (gtx8_txoutclk_i),
        .GTX8_TXRESET_IN                (!ck_160_plllkdet),
        .GTX8_TXUSRCLK2_IN              (snap_clk2),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GTX8_TXN_OUT                   (TXN[3]),
        .GTX8_TXP_OUT                   (TXP[3]),
        .gtx8_force_error               (force_err_wait & force_err_flag[3]),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .GTX8_TXDLYALIGNDISABLE_IN      (gtx8_txdlyaligndisable_i),
        .GTX8_TXDLYALIGNMONENB_IN       (gtx8_txdlyalignmonenb_i),
        .GTX8_TXDLYALIGNMONITOR_OUT     (gtx8_txdlyalignmonitor_i),
        .GTX8_TXDLYALIGNRESET_IN        (gtx8_txdlyalignreset_i),
        .GTX8_TXENPMAPHASEALIGN_IN      (gtx8_txenpmaphasealign_i),
        .GTX8_TXPMASETPHASE_IN          (gtx8_txpmasetphase_i),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTX8_GTXTXRESET_IN             (gtx8_gtxtxreset_i),
        .GTX8_TXRESETDONE_OUT           (gtx8_txresetdone_i),


 
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GTX9  (X0Y9)
        //---------------------- Loopback and Powerdown Ports ----------------------
//jg        .GTX9_RXPOWERDOWN_IN            (gtx9_rxpowerdown_i),
//jg        .GTX9_TXPOWERDOWN_IN            (gtx9_txpowerdown_i),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .GTX9_RXCLKCORCNT_OUT           (gtx9_rxclkcorcnt_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .GTX9_RXBYTEREALIGN_OUT         (gtx9_rxbyterealign_i),
        .GTX9_RXCOMMADET_OUT            (gtx9_rxcommadet_i),
        .GTX9_RXENMCOMMAALIGN_IN        (snap_commaalign),
        .GTX9_RXENPCOMMAALIGN_IN        (snap_commaalign),
        //----------------- Receive Ports - RX Data Path interface -----------------
//jg        .GTX9_RXDATA_OUT                (gtx9_rxdata_i),
        .GTX9_RXRESET_IN                (!ck_160_plllkdet),
        .GTX9_RXUSRCLK2_IN              (snap_clk2),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .GTX9_RXCDRRESET_IN             (gtx9_rxcdrreset_i),
        .GTX9_RXN_IN                    (RXN[5]),
        .GTX9_RXP_IN                    (RXP[5]),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .GTX9_RXLOSSOFSYNC_OUT          (gtx9_rxlossofsync_i),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTX9_GTXRXRESET_IN             (gtx9_gtxrxreset_i),
        .GTX9_MGTREFCLKRX_IN            (q1_clk1_refclk_i),
        .GTX9_PLLRXRESET_IN             (gtx9_pllrxreset_i),
        .GTX9_RXPLLLKDET_OUT            (gtx9_rxplllkdet_i),
        .GTX9_RXRESETDONE_OUT           (gtx9_rxresetdone_i),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .GTX9_RXVALID_OUT               (gtx9_rxvalid_i),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .GTX9_RXPOLARITY_IN             (gtx9_rxpolarity_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GTX9_SEED_IN                 (seed_in[4]),
        .GTX9_RXSEED                  (seed_in[5]),
        .GTX9_TXOUTCLK_OUT              (gtx9_txoutclk_i),
        .GTX9_TXRESET_IN                (!ck_160_plllkdet),
        .GTX9_TXUSRCLK2_IN              (snap_clk2),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GTX9_TXN_OUT                   (TXN[4]),
        .GTX9_TXP_OUT                   (TXP[4]),
        .gtx9_force_error               (force_err_wait & force_err_flag[4]),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .GTX9_TXDLYALIGNDISABLE_IN      (gtx9_txdlyaligndisable_i),
        .GTX9_TXDLYALIGNMONENB_IN       (gtx9_txdlyalignmonenb_i),
        .GTX9_TXDLYALIGNMONITOR_OUT     (gtx9_txdlyalignmonitor_i),
        .GTX9_TXDLYALIGNRESET_IN        (gtx9_txdlyalignreset_i),
        .GTX9_TXENPMAPHASEALIGN_IN      (gtx9_txenpmaphasealign_i),
        .GTX9_TXPMASETPHASE_IN          (gtx9_txpmasetphase_i),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTX9_GTXTXRESET_IN             (gtx9_gtxtxreset_i),
        .GTX9_TXRESETDONE_OUT           (gtx9_txresetdone_i),


 
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GTX10  (X0Y10)
        //---------------------- Loopback and Powerdown Ports ----------------------
//jg        .GTX10_RXPOWERDOWN_IN           (gtx10_rxpowerdown_i),
//jg        .GTX10_TXPOWERDOWN_IN           (gtx10_txpowerdown_i),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .GTX10_RXCLKCORCNT_OUT          (gtx10_rxclkcorcnt_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .GTX10_RXBYTEREALIGN_OUT        (gtx10_rxbyterealign_i),
        .GTX10_RXCOMMADET_OUT           (gtx10_rxcommadet_i),
        .GTX10_RXENMCOMMAALIGN_IN       (snap_commaalign),
        .GTX10_RXENPCOMMAALIGN_IN       (snap_commaalign),
        //----------------- Receive Ports - RX Data Path interface -----------------
//jg        .GTX10_RXDATA_OUT               (gtx10_rxdata_i),
        .GTX10_RXRESET_IN               (!ck_160_plllkdet),
        .GTX10_RXUSRCLK2_IN             (snap_clk2),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .GTX10_RXCDRRESET_IN            (gtx10_rxcdrreset_i),
        .GTX10_RXN_IN                   (RXN[6]),
        .GTX10_RXP_IN                   (RXP[6]),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .GTX10_RXLOSSOFSYNC_OUT         (gtx10_rxlossofsync_i),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTX10_GTXRXRESET_IN            (gtx10_gtxrxreset_i),
        .GTX10_MGTREFCLKRX_IN           (q1_clk1_refclk_i),
        .GTX10_PLLRXRESET_IN            (gtx10_pllrxreset_i),
        .GTX10_RXPLLLKDET_OUT           (gtx10_rxplllkdet_i),
        .GTX10_RXRESETDONE_OUT          (gtx10_rxresetdone_i),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .GTX10_RXVALID_OUT              (gtx10_rxvalid_i),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .GTX10_RXPOLARITY_IN            (gtx10_rxpolarity_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GTX10_SEED_IN                 (seed_in[5]),
        .GTX10_RXSEED                  (seed_in[6]),
        .GTX10_TXOUTCLK_OUT             (gtx10_txoutclk_i),
        .GTX10_TXRESET_IN               (!ck_160_plllkdet),
        .GTX10_TXUSRCLK2_IN             (snap_clk2),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GTX10_TXN_OUT                  (TXN[5]),
        .GTX10_TXP_OUT                  (TXP[5]),
        .gtx10_force_error              (force_err_wait & force_err_flag[5]),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .GTX10_TXDLYALIGNDISABLE_IN     (gtx10_txdlyaligndisable_i),
        .GTX10_TXDLYALIGNMONENB_IN      (gtx10_txdlyalignmonenb_i),
        .GTX10_TXDLYALIGNMONITOR_OUT    (gtx10_txdlyalignmonitor_i),
        .GTX10_TXDLYALIGNRESET_IN       (gtx10_txdlyalignreset_i),
        .GTX10_TXENPMAPHASEALIGN_IN     (gtx10_txenpmaphasealign_i),
        .GTX10_TXPMASETPHASE_IN         (gtx10_txpmasetphase_i),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTX10_GTXTXRESET_IN            (gtx10_gtxtxreset_i),
        .GTX10_TXRESETDONE_OUT          (gtx10_txresetdone_i),


 
 
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GTX11  (X0Y11)
        //---------------------- Loopback and Powerdown Ports ----------------------
//jg        .GTX11_RXPOWERDOWN_IN           (gtx11_rxpowerdown_i),
//jg        .GTX11_TXPOWERDOWN_IN           (gtx11_txpowerdown_i),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .GTX11_RXCLKCORCNT_OUT          (gtx11_rxclkcorcnt_i),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .GTX11_RXBYTEREALIGN_OUT        (gtx11_rxbyterealign_i),
        .GTX11_RXCOMMADET_OUT           (gtx11_rxcommadet_i),
        .GTX11_RXENMCOMMAALIGN_IN       (snap_commaalign),
        .GTX11_RXENPCOMMAALIGN_IN       (snap_commaalign),
        //----------------- Receive Ports - RX Data Path interface -----------------
//jg        .GTX11_RXDATA_OUT               (gtx11_rxdata_i),
        .GTX11_RXRESET_IN               (!ck_160_plllkdet),
        .GTX11_RXUSRCLK2_IN             (snap_clk2),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .GTX11_RXCDRRESET_IN            (gtx11_rxcdrreset_i),
        .GTX11_RXN_IN                   (RXN[7]),
        .GTX11_RXP_IN                   (RXP[7]),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .GTX11_RXLOSSOFSYNC_OUT         (gtx11_rxlossofsync_i),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTX11_GTXRXRESET_IN            (gtx11_gtxrxreset_i),
        .GTX11_MGTREFCLKRX_IN           (q1_clk1_refclk_i),
        .GTX11_PLLRXRESET_IN            (gtx11_pllrxreset_i),
        .GTX11_RXPLLLKDET_OUT           (gtx11_rxplllkdet_i),
        .GTX11_RXRESETDONE_OUT          (gtx11_rxresetdone_i),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .GTX11_RXVALID_OUT              (gtx11_rxvalid_i),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .GTX11_RXPOLARITY_IN            (gtx11_rxpolarity_i),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GTX11_SEED_IN                 (seed_in[6]),
        .GTX11_RXSEED                  (seed_in[7]),
        .GTX11_TXOUTCLK_OUT             (gtx11_txoutclk_i),
        .GTX11_TXRESET_IN               (!ck_160_plllkdet),
        .GTX11_TXUSRCLK2_IN             (snap_clk2),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GTX11_TXN_OUT                  (TXN[6]),
        .GTX11_TXP_OUT                  (TXP[6]),
        .gtx11_force_error              (force_err_wait & force_err_flag[6]),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .GTX11_TXDLYALIGNDISABLE_IN     (gtx11_txdlyaligndisable_i),
        .GTX11_TXDLYALIGNMONENB_IN      (gtx11_txdlyalignmonenb_i),
        .GTX11_TXDLYALIGNMONITOR_OUT    (gtx11_txdlyalignmonitor_i),
        .GTX11_TXDLYALIGNRESET_IN       (gtx11_txdlyalignreset_i),
        .GTX11_TXENPMAPHASEALIGN_IN     (gtx11_txenpmaphasealign_i),
        .GTX11_TXPMASETPHASE_IN         (gtx11_txpmasetphase_i),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTX11_GTXTXRESET_IN            (gtx11_gtxtxreset_i),
        .GTX11_TXRESETDONE_OUT          (gtx11_txresetdone_i)


    );


    //---------------------------- TXSYNC module ------------------------------
    // The TXSYNC module performs phase synchronization for all the active TX datapaths. It
    // waits for the user clocks to be stable, then drives the phase align signals on each
    // GTX. When phase synchronization is complete, it asserts SYNC_DONE
    
    // Include the TX_SYNC module in your own design to perform phase synchronization if
    // your protocol bypasses the TX Buffers
  

    // SIM_TXPMASETPHASE_SPEEDUP is a simulation only attribute and MUST be set to 0 
    // during implementation     
    TX_SYNC #
    (
        .SIM_TXPMASETPHASE_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP)
    )
    gtx0_txsync_i 
    (
        .TXENPMAPHASEALIGN(gtx0_txenpmaphasealign_i), // OUT to GTX
        .TXPMASETPHASE(gtx0_txpmasetphase_i),         // OUT to GTX
        .TXDLYALIGNDISABLE(gtx0_txdlyaligndisable_i), // OUT to GTX
        .TXDLYALIGNRESET(gtx0_txdlyalignreset_i),     // OUT to GTX
        .SYNC_DONE(gtx0_tx_sync_done_i),              // OUT to reset "data transmit logic"
        .USER_CLK(snap_clk2),                         // input
        .RESET(!gtx0_txresetdone_r2)                  // input
    );


    // SIM_TXPMASETPHASE_SPEEDUP is a simulation only attribute and MUST be set to 0 
    // during implementation     
    TX_SYNC #
    (
        .SIM_TXPMASETPHASE_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP)
    )
    gtx1_txsync_i 
    (
        .TXENPMAPHASEALIGN(gtx1_txenpmaphasealign_i),
        .TXPMASETPHASE(gtx1_txpmasetphase_i),
        .TXDLYALIGNDISABLE(gtx1_txdlyaligndisable_i),
        .TXDLYALIGNRESET(gtx1_txdlyalignreset_i),
        .SYNC_DONE(gtx1_tx_sync_done_i),
        .USER_CLK(snap_clk2),
        .RESET(!gtx1_txresetdone_r2)
    );


    // SIM_TXPMASETPHASE_SPEEDUP is a simulation only attribute and MUST be set to 0 
    // during implementation     
    TX_SYNC #
    (
        .SIM_TXPMASETPHASE_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP)
    )
    gtx2_txsync_i 
    (
        .TXENPMAPHASEALIGN(gtx2_txenpmaphasealign_i),
        .TXPMASETPHASE(gtx2_txpmasetphase_i),
        .TXDLYALIGNDISABLE(gtx2_txdlyaligndisable_i),
        .TXDLYALIGNRESET(gtx2_txdlyalignreset_i),
        .SYNC_DONE(syncdone_snapt[7]),
        .USER_CLK(snap_clk2),
        .RESET(!gtx2_txresetdone_r2)
    );


    // SIM_TXPMASETPHASE_SPEEDUP is a simulation only attribute and MUST be set to 0 
    // during implementation     
    TX_SYNC #
    (
        .SIM_TXPMASETPHASE_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP)
    )
    gtx3_txsync_i 
    (
        .TXENPMAPHASEALIGN(gtx3_txenpmaphasealign_i),
        .TXPMASETPHASE(gtx3_txpmasetphase_i),
        .TXDLYALIGNDISABLE(gtx3_txdlyaligndisable_i),
        .TXDLYALIGNRESET(gtx3_txdlyalignreset_i),
        .SYNC_DONE(syncdone_snapt[0]),
        .USER_CLK(snap_clk2),
        .RESET(!gtx3_txresetdone_r2)
    );


    // SIM_TXPMASETPHASE_SPEEDUP is a simulation only attribute and MUST be set to 0 
    // during implementation     
    TX_SYNC #
    (
        .SIM_TXPMASETPHASE_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP)
    )
    gtx4_txsync_i 
    (
        .TXENPMAPHASEALIGN(gtx4_txenpmaphasealign_i),
        .TXPMASETPHASE(gtx4_txpmasetphase_i),
        .TXDLYALIGNDISABLE(gtx4_txdlyaligndisable_i),
        .TXDLYALIGNRESET(gtx4_txdlyalignreset_i),
        .SYNC_DONE(syncdone_snapt[1]),
        .USER_CLK(snap_clk2),
        .RESET(!gtx4_txresetdone_r2)
    );


    // SIM_TXPMASETPHASE_SPEEDUP is a simulation only attribute and MUST be set to 0 
    // during implementation     
    TX_SYNC #
    (
        .SIM_TXPMASETPHASE_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP)
    )
    gtx5_txsync_i 
    (
        .TXENPMAPHASEALIGN(gtx5_txenpmaphasealign_i),
        .TXPMASETPHASE(gtx5_txpmasetphase_i),
        .TXDLYALIGNDISABLE(gtx5_txdlyaligndisable_i),
        .TXDLYALIGNRESET(gtx5_txdlyalignreset_i),
        .SYNC_DONE(gtx5_tx_sync_done_i),
        .USER_CLK(snap_clk2),
        .RESET(!gtx5_txresetdone_r2)
    );


    // SIM_TXPMASETPHASE_SPEEDUP is a simulation only attribute and MUST be set to 0 
    // during implementation     
    TX_SYNC #
    (
        .SIM_TXPMASETPHASE_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP)
    )
    gtx6_txsync_i 
    (
        .TXENPMAPHASEALIGN(gtx6_txenpmaphasealign_i),
        .TXPMASETPHASE(gtx6_txpmasetphase_i),
        .TXDLYALIGNDISABLE(gtx6_txdlyaligndisable_i),
        .TXDLYALIGNRESET(gtx6_txdlyalignreset_i),
        .SYNC_DONE(gtx6_tx_sync_done_i),
        .USER_CLK(snap_clk2),
        .RESET(!gtx6_txresetdone_r2)
    );


    // SIM_TXPMASETPHASE_SPEEDUP is a simulation only attribute and MUST be set to 0 
    // during implementation     
    TX_SYNC #
    (
        .SIM_TXPMASETPHASE_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP)
    )
    gtx7_txsync_i 
    (
        .TXENPMAPHASEALIGN(gtx7_txenpmaphasealign_i),
        .TXPMASETPHASE(gtx7_txpmasetphase_i),
        .TXDLYALIGNDISABLE(gtx7_txdlyaligndisable_i),
        .TXDLYALIGNRESET(gtx7_txdlyalignreset_i),
        .SYNC_DONE(syncdone_snapt[2]),
        .USER_CLK(snap_clk2),
        .RESET(!gtx7_txresetdone_r2)
    );


    // SIM_TXPMASETPHASE_SPEEDUP is a simulation only attribute and MUST be set to 0 
    // during implementation     
    TX_SYNC #
    (
        .SIM_TXPMASETPHASE_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP)
    )
    gtx8_txsync_i 
    (
        .TXENPMAPHASEALIGN(gtx8_txenpmaphasealign_i),
        .TXPMASETPHASE(gtx8_txpmasetphase_i),
        .TXDLYALIGNDISABLE(gtx8_txdlyaligndisable_i),
        .TXDLYALIGNRESET(gtx8_txdlyalignreset_i),
        .SYNC_DONE(syncdone_snapt[3]),
        .USER_CLK(snap_clk2),
        .RESET(!gtx8_txresetdone_r2)
    );


    // SIM_TXPMASETPHASE_SPEEDUP is a simulation only attribute and MUST be set to 0 
    // during implementation     
    TX_SYNC #
    (
        .SIM_TXPMASETPHASE_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP)
    )
    gtx9_txsync_i 
    (
        .TXENPMAPHASEALIGN(gtx9_txenpmaphasealign_i),
        .TXPMASETPHASE(gtx9_txpmasetphase_i),
        .TXDLYALIGNDISABLE(gtx9_txdlyaligndisable_i),
        .TXDLYALIGNRESET(gtx9_txdlyalignreset_i),
        .SYNC_DONE(syncdone_snapt[4]),
        .USER_CLK(snap_clk2),
        .RESET(!gtx9_txresetdone_r2)
    );


    // SIM_TXPMASETPHASE_SPEEDUP is a simulation only attribute and MUST be set to 0 
    // during implementation     
    TX_SYNC #
    (
        .SIM_TXPMASETPHASE_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP)
    )
    gtx10_txsync_i 
    (
        .TXENPMAPHASEALIGN(gtx10_txenpmaphasealign_i),
        .TXPMASETPHASE(gtx10_txpmasetphase_i),
        .TXDLYALIGNDISABLE(gtx10_txdlyaligndisable_i),
        .TXDLYALIGNRESET(gtx10_txdlyalignreset_i),
        .SYNC_DONE(syncdone_snapt[5]),
        .USER_CLK(snap_clk2),
        .RESET(!gtx10_txresetdone_r2)
    );


    // SIM_TXPMASETPHASE_SPEEDUP is a simulation only attribute and MUST be set to 0 
    // during implementation     
    TX_SYNC #
    (
        .SIM_TXPMASETPHASE_SPEEDUP   (EXAMPLE_SIM_GTXRESET_SPEEDUP)
    )
    gtx11_txsync_i 
    (
        .TXENPMAPHASEALIGN(gtx11_txenpmaphasealign_i),
        .TXPMASETPHASE(gtx11_txpmasetphase_i),
        .TXDLYALIGNDISABLE(gtx11_txdlyaligndisable_i),
        .TXDLYALIGNRESET(gtx11_txdlyalignreset_i),
        .SYNC_DONE(syncdone_snapt[6]),
        .USER_CLK(snap_clk2),
        .RESET(!gtx11_txresetdone_r2)
    );

    


    //------------------------ User Module Resets -----------------------------
    // All the User Modules i.e. FRAME_GEN, FRAME_CHECK and the sync modules
    // are held in reset till the RESETDONE goes high. 
    // The RESETDONE is registered a couple of times on *USRCLK2 and connected 
    // to the reset of the modules
    

//jghere
//    assign all_rx_ready = gtx4_rxresetdone_r3 & gtx5_rxresetdone_r3 & gtx6_rxresetdone_r3 & gtx7_rxresetdone_r3 & gtx8_rxresetdone_r3 & gtx9_rxresetdone_r3 & gtx10_rxresetdone_r3 & gtx11_rxresetdone_r3;
    assign all_rx_ready = gtx0_rxresetdone_r3 & gtx1_rxresetdone_r3 & gtx2_rxresetdone_r3 & gtx3_rxresetdone_r3 & gtx8_rxresetdone_r3 & gtx9_rxresetdone_r3 & gtx10_rxresetdone_r3 & gtx11_rxresetdone_r3;
    assign all_tx_ready = gtx3_txresetdone_r2 & gtx4_txresetdone_r2 & gtx7_txresetdone_r2 & gtx8_txresetdone_r2 & gtx9_txresetdone_r2 & gtx10_txresetdone_r2 & gtx11_txresetdone_r2 & gtx2_txresetdone_r2;

    always @(posedge snap_clk2)
            gtx0_rxresetdone_i_r   <=   `DLY gtx0_rxresetdone_i;

    always @(posedge snap_clk2 or negedge gtx0_rxresetdone_i_r)

    begin
        if (!gtx0_rxresetdone_i_r)
        begin
            gtx0_rxresetdone_r      <=   `DLY 1'b0;
            gtx0_rxresetdone_r2     <=   `DLY 1'b0;
        end
        else
        begin
            gtx0_rxresetdone_r      <=   `DLY gtx0_rxresetdone_i_r;
            gtx0_rxresetdone_r2     <=   `DLY gtx0_rxresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx0_rxresetdone_r3   <=   `DLY gtx0_rxresetdone_r2;
    
    
    always @(posedge snap_clk2 or negedge gtx0_txresetdone_i)

    begin
        if (!gtx0_txresetdone_i)
        begin
            gtx0_txresetdone_r    <=   `DLY 1'b0;
            gtx0_txresetdone_r2   <=   `DLY 1'b0;
        end
        else
        begin
            gtx0_txresetdone_r    <=   `DLY gtx0_txresetdone_i;
            gtx0_txresetdone_r2   <=   `DLY gtx0_txresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx1_rxresetdone_i_r   <=   `DLY gtx1_rxresetdone_i;

    always @(posedge snap_clk2 or negedge gtx1_rxresetdone_i_r)

    begin
        if (!gtx1_rxresetdone_i_r)
        begin
            gtx1_rxresetdone_r      <=   `DLY 1'b0;
            gtx1_rxresetdone_r2     <=   `DLY 1'b0;
        end
        else
        begin
            gtx1_rxresetdone_r      <=   `DLY gtx1_rxresetdone_i_r;
            gtx1_rxresetdone_r2     <=   `DLY gtx1_rxresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx1_rxresetdone_r3   <=   `DLY gtx1_rxresetdone_r2;
    
    
    always @(posedge snap_clk2 or negedge gtx1_txresetdone_i)

    begin
        if (!gtx1_txresetdone_i)
        begin
            gtx1_txresetdone_r    <=   `DLY 1'b0;
            gtx1_txresetdone_r2   <=   `DLY 1'b0;
        end
        else
        begin
            gtx1_txresetdone_r    <=   `DLY gtx1_txresetdone_i;
            gtx1_txresetdone_r2   <=   `DLY gtx1_txresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx2_rxresetdone_i_r   <=   `DLY gtx2_rxresetdone_i;

    always @(posedge snap_clk2 or negedge gtx2_rxresetdone_i_r)

    begin
        if (!gtx2_rxresetdone_i_r)
        begin
            gtx2_rxresetdone_r      <=   `DLY 1'b0;
            gtx2_rxresetdone_r2     <=   `DLY 1'b0;
        end
        else
        begin
            gtx2_rxresetdone_r      <=   `DLY gtx2_rxresetdone_i_r;
            gtx2_rxresetdone_r2     <=   `DLY gtx2_rxresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx2_rxresetdone_r3   <=   `DLY gtx2_rxresetdone_r2;
    
    
    always @(posedge snap_clk2 or negedge gtx2_txresetdone_i)

    begin
        if (!gtx2_txresetdone_i)
        begin
            gtx2_txresetdone_r    <=   `DLY 1'b0;
            gtx2_txresetdone_r2   <=   `DLY 1'b0;
        end
        else
        begin
            gtx2_txresetdone_r    <=   `DLY gtx2_txresetdone_i;
            gtx2_txresetdone_r2   <=   `DLY gtx2_txresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx3_rxresetdone_i_r   <=   `DLY gtx3_rxresetdone_i;

    always @(posedge snap_clk2 or negedge gtx3_rxresetdone_i_r)

    begin
        if (!gtx3_rxresetdone_i_r)
        begin
            gtx3_rxresetdone_r      <=   `DLY 1'b0;
            gtx3_rxresetdone_r2     <=   `DLY 1'b0;
        end
        else
        begin
            gtx3_rxresetdone_r      <=   `DLY gtx3_rxresetdone_i_r;
            gtx3_rxresetdone_r2     <=   `DLY gtx3_rxresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx3_rxresetdone_r3   <=   `DLY gtx3_rxresetdone_r2;
    
    
    always @(posedge snap_clk2 or negedge gtx3_txresetdone_i)

    begin
        if (!gtx3_txresetdone_i)
        begin
            gtx3_txresetdone_r    <=   `DLY 1'b0;
            gtx3_txresetdone_r2   <=   `DLY 1'b0;
        end
        else
        begin
            gtx3_txresetdone_r    <=   `DLY gtx3_txresetdone_i;
            gtx3_txresetdone_r2   <=   `DLY gtx3_txresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx4_rxresetdone_i_r   <=   `DLY gtx4_rxresetdone_i;

    always @(posedge snap_clk2 or negedge gtx4_rxresetdone_i_r)

    begin
        if (!gtx4_rxresetdone_i_r)
        begin
            gtx4_rxresetdone_r      <=   `DLY 1'b0;
            gtx4_rxresetdone_r2     <=   `DLY 1'b0;
        end
        else
        begin
            gtx4_rxresetdone_r      <=   `DLY gtx4_rxresetdone_i_r;
            gtx4_rxresetdone_r2     <=   `DLY gtx4_rxresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx4_rxresetdone_r3   <=   `DLY gtx4_rxresetdone_r2;
    
    
    always @(posedge snap_clk2 or negedge gtx4_txresetdone_i)

    begin
        if (!gtx4_txresetdone_i)
        begin
            gtx4_txresetdone_r    <=   `DLY 1'b0;
            gtx4_txresetdone_r2   <=   `DLY 1'b0;
        end
        else
        begin
            gtx4_txresetdone_r    <=   `DLY gtx4_txresetdone_i;
            gtx4_txresetdone_r2   <=   `DLY gtx4_txresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx5_rxresetdone_i_r   <=   `DLY gtx5_rxresetdone_i;

    always @(posedge snap_clk2 or negedge gtx5_rxresetdone_i_r)

    begin
        if (!gtx5_rxresetdone_i_r)
        begin
            gtx5_rxresetdone_r      <=   `DLY 1'b0;
            gtx5_rxresetdone_r2     <=   `DLY 1'b0;
        end
        else
        begin
            gtx5_rxresetdone_r      <=   `DLY gtx5_rxresetdone_i_r;
            gtx5_rxresetdone_r2     <=   `DLY gtx5_rxresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx5_rxresetdone_r3   <=   `DLY gtx5_rxresetdone_r2;
    
    
    always @(posedge snap_clk2 or negedge gtx5_txresetdone_i)

    begin
        if (!gtx5_txresetdone_i)
        begin
            gtx5_txresetdone_r    <=   `DLY 1'b0;
            gtx5_txresetdone_r2   <=   `DLY 1'b0;
        end
        else
        begin
            gtx5_txresetdone_r    <=   `DLY gtx5_txresetdone_i;
            gtx5_txresetdone_r2   <=   `DLY gtx5_txresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx6_rxresetdone_i_r   <=   `DLY gtx6_rxresetdone_i;

    always @(posedge snap_clk2 or negedge gtx6_rxresetdone_i_r)

    begin
        if (!gtx6_rxresetdone_i_r)
        begin
            gtx6_rxresetdone_r      <=   `DLY 1'b0;
            gtx6_rxresetdone_r2     <=   `DLY 1'b0;
        end
        else
        begin
            gtx6_rxresetdone_r      <=   `DLY gtx6_rxresetdone_i_r;
            gtx6_rxresetdone_r2     <=   `DLY gtx6_rxresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx6_rxresetdone_r3   <=   `DLY gtx6_rxresetdone_r2;
    
    
    always @(posedge snap_clk2 or negedge gtx6_txresetdone_i)

    begin
        if (!gtx6_txresetdone_i)
        begin
            gtx6_txresetdone_r    <=   `DLY 1'b0;
            gtx6_txresetdone_r2   <=   `DLY 1'b0;
        end
        else
        begin
            gtx6_txresetdone_r    <=   `DLY gtx6_txresetdone_i;
            gtx6_txresetdone_r2   <=   `DLY gtx6_txresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx7_rxresetdone_i_r   <=   `DLY gtx7_rxresetdone_i;

    always @(posedge snap_clk2 or negedge gtx7_rxresetdone_i_r)

    begin
        if (!gtx7_rxresetdone_i_r)
        begin
            gtx7_rxresetdone_r      <=   `DLY 1'b0;
            gtx7_rxresetdone_r2     <=   `DLY 1'b0;
        end
        else
        begin
            gtx7_rxresetdone_r      <=   `DLY gtx7_rxresetdone_i_r;
            gtx7_rxresetdone_r2     <=   `DLY gtx7_rxresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx7_rxresetdone_r3   <=   `DLY gtx7_rxresetdone_r2;
    
    
    always @(posedge snap_clk2 or negedge gtx7_txresetdone_i)

    begin
        if (!gtx7_txresetdone_i)
        begin
            gtx7_txresetdone_r    <=   `DLY 1'b0;
            gtx7_txresetdone_r2   <=   `DLY 1'b0;
        end
        else
        begin
            gtx7_txresetdone_r    <=   `DLY gtx7_txresetdone_i;
            gtx7_txresetdone_r2   <=   `DLY gtx7_txresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx8_rxresetdone_i_r   <=   `DLY gtx8_rxresetdone_i;

    always @(posedge snap_clk2 or negedge gtx8_rxresetdone_i_r)

    begin
        if (!gtx8_rxresetdone_i_r)
        begin
            gtx8_rxresetdone_r      <=   `DLY 1'b0;
            gtx8_rxresetdone_r2     <=   `DLY 1'b0;
        end
        else
        begin
            gtx8_rxresetdone_r      <=   `DLY gtx8_rxresetdone_i_r;
            gtx8_rxresetdone_r2     <=   `DLY gtx8_rxresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx8_rxresetdone_r3   <=   `DLY gtx8_rxresetdone_r2;
    
    
    always @(posedge snap_clk2 or negedge gtx8_txresetdone_i)

    begin
        if (!gtx8_txresetdone_i)
        begin
            gtx8_txresetdone_r    <=   `DLY 1'b0;
            gtx8_txresetdone_r2   <=   `DLY 1'b0;
        end
        else
        begin
            gtx8_txresetdone_r    <=   `DLY gtx8_txresetdone_i;
            gtx8_txresetdone_r2   <=   `DLY gtx8_txresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx9_rxresetdone_i_r   <=   `DLY gtx9_rxresetdone_i;

    always @(posedge snap_clk2 or negedge gtx9_rxresetdone_i_r)

    begin
        if (!gtx9_rxresetdone_i_r)
        begin
            gtx9_rxresetdone_r      <=   `DLY 1'b0;
            gtx9_rxresetdone_r2     <=   `DLY 1'b0;
        end
        else
        begin
            gtx9_rxresetdone_r      <=   `DLY gtx9_rxresetdone_i_r;
            gtx9_rxresetdone_r2     <=   `DLY gtx9_rxresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx9_rxresetdone_r3   <=   `DLY gtx9_rxresetdone_r2;
    
    
    always @(posedge snap_clk2 or negedge gtx9_txresetdone_i)

    begin
        if (!gtx9_txresetdone_i)
        begin
            gtx9_txresetdone_r    <=   `DLY 1'b0;
            gtx9_txresetdone_r2   <=   `DLY 1'b0;
        end
        else
        begin
            gtx9_txresetdone_r    <=   `DLY gtx9_txresetdone_i;
            gtx9_txresetdone_r2   <=   `DLY gtx9_txresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx10_rxresetdone_i_r   <=   `DLY gtx10_rxresetdone_i;

    always @(posedge snap_clk2 or negedge gtx10_rxresetdone_i_r)

    begin
        if (!gtx10_rxresetdone_i_r)
        begin
            gtx10_rxresetdone_r      <=   `DLY 1'b0;
            gtx10_rxresetdone_r2     <=   `DLY 1'b0;
        end
        else
        begin
            gtx10_rxresetdone_r      <=   `DLY gtx10_rxresetdone_i_r;
            gtx10_rxresetdone_r2     <=   `DLY gtx10_rxresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx10_rxresetdone_r3   <=   `DLY gtx10_rxresetdone_r2;
    
    
    always @(posedge snap_clk2 or negedge gtx10_txresetdone_i)

    begin
        if (!gtx10_txresetdone_i)
        begin
            gtx10_txresetdone_r    <=   `DLY 1'b0;
            gtx10_txresetdone_r2   <=   `DLY 1'b0;
        end
        else
        begin
            gtx10_txresetdone_r    <=   `DLY gtx10_txresetdone_i;
            gtx10_txresetdone_r2   <=   `DLY gtx10_txresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx11_rxresetdone_i_r   <=   `DLY gtx11_rxresetdone_i;

    always @(posedge snap_clk2 or negedge gtx11_rxresetdone_i_r)

    begin
        if (!gtx11_rxresetdone_i_r)
        begin
            gtx11_rxresetdone_r      <=   `DLY 1'b0;
            gtx11_rxresetdone_r2     <=   `DLY 1'b0;
        end
        else
        begin
            gtx11_rxresetdone_r      <=   `DLY gtx11_rxresetdone_i_r;
            gtx11_rxresetdone_r2     <=   `DLY gtx11_rxresetdone_r;
        end
    end

    always @(posedge snap_clk2)
            gtx11_rxresetdone_r3   <=   `DLY gtx11_rxresetdone_r2;
    
    
    always @(posedge snap_clk2 or negedge gtx11_txresetdone_i)

    begin
        if (!gtx11_txresetdone_i)
        begin
            gtx11_txresetdone_r    <=   `DLY 1'b0;
            gtx11_txresetdone_r2   <=   `DLY 1'b0;
        end
        else
        begin
            gtx11_txresetdone_r    <=   `DLY gtx11_txresetdone_i;
            gtx11_txresetdone_r2   <=   `DLY gtx11_txresetdone_r;
        end
    end


generate
begin: no_chipscope

    // If Chipscope is not being used, drive GTX reset signal
    // from the top level ports
    assign  gtx0_gtxrxreset_i = GTXRXRESET_IN;
    assign  gtx0_gtxtxreset_i = GTXTXRESET_IN;
    assign  gtx1_gtxrxreset_i = GTXRXRESET_IN;
    assign  gtx1_gtxtxreset_i = GTXTXRESET_IN;
    assign  gtx2_gtxrxreset_i = GTXRXRESET_IN;
    assign  gtx2_gtxtxreset_i = GTXTXRESET_IN;
    assign  gtx3_gtxrxreset_i = GTXRXRESET_IN;
    assign  gtx3_gtxtxreset_i = GTXTXRESET_IN;
    assign  gtx4_gtxrxreset_i = GTXRXRESET_IN;
    assign  gtx4_gtxtxreset_i = GTXTXRESET_IN;
    assign  gtx5_gtxrxreset_i = GTXRXRESET_IN;
    assign  gtx5_gtxtxreset_i = GTXTXRESET_IN;
    assign  gtx6_gtxrxreset_i = GTXRXRESET_IN;
    assign  gtx6_gtxtxreset_i = GTXTXRESET_IN;
    assign  gtx7_gtxrxreset_i = GTXRXRESET_IN;
    assign  gtx7_gtxtxreset_i = GTXTXRESET_IN;
    assign  gtx8_gtxrxreset_i = GTXRXRESET_IN;
    assign  gtx8_gtxtxreset_i = GTXTXRESET_IN;
    assign  gtx9_gtxrxreset_i = GTXRXRESET_IN;
    assign  gtx9_gtxtxreset_i = GTXTXRESET_IN;
    assign  gtx10_gtxrxreset_i = GTXRXRESET_IN;
    assign  gtx10_gtxtxreset_i = GTXTXRESET_IN;
    assign  gtx11_gtxrxreset_i = GTXRXRESET_IN;
    assign  gtx11_gtxtxreset_i = GTXTXRESET_IN;

    // assign resets for frame_check modules
    assign  gtx0_rx_system_reset_c = !gtx0_rxresetdone_r3;
    assign  gtx1_rx_system_reset_c = !gtx1_rxresetdone_r3;
    assign  gtx2_rx_system_reset_c = !gtx2_rxresetdone_r3;
    assign  gtx3_rx_system_reset_c = !gtx3_rxresetdone_r3;
    assign  gtx4_rx_system_reset_c = !gtx4_rxresetdone_r3;
    assign  gtx5_rx_system_reset_c = !gtx5_rxresetdone_r3;
    assign  gtx6_rx_system_reset_c = !gtx6_rxresetdone_r3;
    assign  gtx7_rx_system_reset_c = !gtx7_rxresetdone_r3;
    assign  gtx8_rx_system_reset_c = !gtx8_rxresetdone_r3;
    assign  gtx9_rx_system_reset_c = !gtx9_rxresetdone_r3;
    assign  gtx10_rx_system_reset_c = !gtx10_rxresetdone_r3;
    assign  gtx11_rx_system_reset_c = !gtx11_rxresetdone_r3;

    assign  gtxtxreset_i                         =  tied_to_ground_i;
    assign  gtxrxreset_i                         =  tied_to_ground_i;
    assign  user_tx_reset_i                      =  tied_to_ground_i;
    assign  user_rx_reset_i                      =  tied_to_ground_i;
    assign  mux_sel_i                            =  tied_to_ground_vec_i[3:0];
    assign  gtx0_txdlyalignmonenb_i              =  tied_to_ground_i;
    assign  gtx0_txpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx0_pllrxreset_i                    =  tied_to_ground_i;
    assign  gtx0_rxpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx0_rxcdrreset_i                    =  tied_to_ground_i;
    assign  gtx0_rxpolarity_i                    =  tied_to_ground_i;
    assign  gtx1_txdlyalignmonenb_i              =  tied_to_ground_i;
    assign  gtx1_txpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx1_pllrxreset_i                    =  tied_to_ground_i;
    assign  gtx1_rxpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx1_rxcdrreset_i                    =  tied_to_ground_i;
    assign  gtx1_rxpolarity_i                    =  tied_to_ground_i;
    assign  gtx2_txdlyalignmonenb_i              =  tied_to_ground_i;
    assign  gtx2_txpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx2_pllrxreset_i                    =  tied_to_ground_i;
    assign  gtx2_rxpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx2_rxcdrreset_i                    =  tied_to_ground_i;
    assign  gtx2_rxpolarity_i                    =  tied_to_ground_i;
    assign  gtx3_txdlyalignmonenb_i              =  tied_to_ground_i;
    assign  gtx3_txpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx3_pllrxreset_i                    =  tied_to_ground_i;
    assign  gtx3_rxpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx3_rxcdrreset_i                    =  tied_to_ground_i;
    assign  gtx3_rxpolarity_i                    =  tied_to_ground_i;
    assign  gtx4_txdlyalignmonenb_i              =  tied_to_ground_i;
    assign  gtx4_txpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx4_pllrxreset_i                    =  tied_to_ground_i;
    assign  gtx4_rxpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx4_rxcdrreset_i                    =  tied_to_ground_i;
    assign  gtx4_rxpolarity_i                    =  tied_to_ground_i;
    assign  gtx5_txdlyalignmonenb_i              =  tied_to_ground_i;
    assign  gtx5_txpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx5_pllrxreset_i                    =  tied_to_ground_i;
    assign  gtx5_rxpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx5_rxcdrreset_i                    =  tied_to_ground_i;
    assign  gtx5_rxpolarity_i                    =  tied_to_ground_i;
    assign  gtx6_txdlyalignmonenb_i              =  tied_to_ground_i;
    assign  gtx6_txpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx6_pllrxreset_i                    =  tied_to_ground_i;
    assign  gtx6_rxpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx6_rxcdrreset_i                    =  tied_to_ground_i;
    assign  gtx6_rxpolarity_i                    =  tied_to_ground_i;
    assign  gtx7_txdlyalignmonenb_i              =  tied_to_ground_i;
    assign  gtx7_txpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx7_pllrxreset_i                    =  tied_to_ground_i;
    assign  gtx7_rxpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx7_rxcdrreset_i                    =  tied_to_ground_i;
    assign  gtx7_rxpolarity_i                    =  tied_to_ground_i;
    assign  gtx8_txdlyalignmonenb_i              =  tied_to_ground_i;
    assign  gtx8_txpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx8_pllrxreset_i                    =  tied_to_ground_i;
    assign  gtx8_rxpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx8_rxcdrreset_i                    =  tied_to_ground_i;
    assign  gtx8_rxpolarity_i                    =  tied_to_ground_i;
    assign  gtx9_txdlyalignmonenb_i              =  tied_to_ground_i;
    assign  gtx9_txpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx9_pllrxreset_i                    =  tied_to_ground_i;
    assign  gtx9_rxpowerdown_i                   =  tied_to_ground_vec_i[1:0];
    assign  gtx9_rxcdrreset_i                    =  tied_to_ground_i;
    assign  gtx9_rxpolarity_i                    =  1'b1; // tied_to_ground_i;
    assign  gtx10_txdlyalignmonenb_i             =  tied_to_ground_i;
    assign  gtx10_txpowerdown_i                  =  tied_to_ground_vec_i[1:0];
    assign  gtx10_pllrxreset_i                   =  tied_to_ground_i;
    assign  gtx10_rxpowerdown_i                  =  tied_to_ground_vec_i[1:0];
    assign  gtx10_rxcdrreset_i                   =  tied_to_ground_i;
    assign  gtx10_rxpolarity_i                   =  1'b1; // tied_to_ground_i;
    assign  gtx11_txdlyalignmonenb_i             =  tied_to_ground_i;
    assign  gtx11_txpowerdown_i                  =  tied_to_ground_vec_i[1:0];
    assign  gtx11_pllrxreset_i                   =  tied_to_ground_i;
    assign  gtx11_rxpowerdown_i                  =  tied_to_ground_vec_i[1:0];
    assign  gtx11_rxcdrreset_i                   =  tied_to_ground_i;
    assign  gtx11_rxpolarity_i                   =  tied_to_ground_i;


end
endgenerate //End generate for EXAMPLE_USE_CHIPSCOPE


endmodule

