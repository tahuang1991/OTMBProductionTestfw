------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 1.8
--  \   \         Application : Virtex-6 FPGA GTX Transceiver Wizard 
--  /   /         Filename : trg_tx_buf_bypass_top.vhd
-- /___/   /\     Timestamp : 
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module TRG_TX_BUF_BYPASS_TOP
-- Generated by Xilinx Virtex-6 FPGA GTX Transceiver Wizard
-- 
-- 
-- (c) Copyright 2009-2010 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***********************************Entity Declaration************************

entity TRG_TX_BUF_BYPASS_TOP is
generic
(
    EXAMPLE_CONFIG_INDEPENDENT_LANES        : integer   := 1;
    EXAMPLE_LANE_WITH_START_CHAR            : integer   := 0;    -- specifies lane with unique start frame ch
    EXAMPLE_WORDS_IN_BRAM                   : integer   := 512;  -- specifies amount of data in BRAM
    EXAMPLE_SIM_GTXRESET_SPEEDUP            : integer   := 0;    -- simulation setting for GTX SecureIP model
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 1     -- Set to 1 to use Chipscope to drive resets
);
port
(
    Q1_CLK1_MGTREFCLK_PAD_N_IN              : in   std_logic;
    Q1_CLK1_MGTREFCLK_PAD_P_IN              : in   std_logic;
    GTXTXRESET_IN                           : in   std_logic;
    GTXRXRESET_IN                           : in   std_logic;
    RXN_IN                                  : in   std_logic;
    RXP_IN                                  : in   std_logic;
    TXN_OUT                                 : out  std_logic;
    TXP_OUT                                 : out  std_logic
    
);


end TRG_TX_BUF_BYPASS_TOP;
    
architecture RTL of TRG_TX_BUF_BYPASS_TOP is

--**************************Component Declarations*****************************


component TRG_TX_BUF_BYPASS 
generic
(
    -- Simulation attributes
    WRAPPER_SIM_GTXRESET_SPEEDUP    : integer   := 0 -- Set to 1 to speed up sim reset
);
port
(

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GTX0  (X0_Y2)

    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    GTX0_RXN_IN                             : in   std_logic;
    GTX0_RXP_IN                             : in   std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    GTX0_TXCHARISK_IN                       : in   std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GTX0_TXDATA_IN                          : in   std_logic_vector(31 downto 0);
    GTX0_TXOUTCLK_OUT                       : out  std_logic;
    GTX0_TXUSRCLK_IN                        : in   std_logic;
    GTX0_TXUSRCLK2_IN                       : in   std_logic;
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GTX0_TXN_OUT                            : out  std_logic;
    GTX0_TXP_OUT                            : out  std_logic;
    -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    GTX0_TXDLYALIGNDISABLE_IN               : in   std_logic;
    GTX0_TXDLYALIGNMONENB_IN                : in   std_logic;
    GTX0_TXDLYALIGNMONITOR_OUT              : out  std_logic_vector(7 downto 0);
    GTX0_TXDLYALIGNRESET_IN                 : in   std_logic;
    GTX0_TXENPMAPHASEALIGN_IN               : in   std_logic;
    GTX0_TXPMASETPHASE_IN                   : in   std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    GTX0_GTXTXRESET_IN                      : in   std_logic;
    GTX0_MGTREFCLKTX_IN                     : in   std_logic;
    GTX0_PLLTXRESET_IN                      : in   std_logic;
    GTX0_TXPLLLKDET_OUT                     : out  std_logic;
    GTX0_TXRESETDONE_OUT                    : out  std_logic


);
end component;

component MGT_USRCLK_SOURCE 
generic
(
    FREQUENCY_MODE   : string   := "LOW";    
    PERFORMANCE_MODE : string   := "MAX_SPEED"    
);
port
(
    DIV1_OUT                : out std_logic;
    DIV2_OUT                : out std_logic;
    DCM_LOCKED_OUT          : out std_logic;
    CLK_IN                  : in  std_logic;
    DCM_RESET_IN            : in  std_logic

);
end component;

component FRAME_GEN 
generic
(
    WORDS_IN_BRAM : integer    :=   256;
    MEM_00       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_01       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_02       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_03       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_04       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_05       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_06       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_07       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_08       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_09       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_10       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_11       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_12       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_13       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_14       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_15       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_16       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_17       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_18       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_19       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_20       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_21       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_22       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_23       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_24       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_25       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_26       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_27       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_28       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_29       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_30       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_31       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_32       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_33       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_34       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_35       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_36       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_37       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_38       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_39       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_00      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_01      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_02      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_03      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_04      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_05      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_06      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_07      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000"
);    
port
(
    -- User Interface
    TX_DATA             : out   std_logic_vector(39 downto 0);
    TX_CHARISK          : out   std_logic_vector(3 downto 0); 

    -- System Interface
    USER_CLK            : in    std_logic;
    SYSTEM_RESET        : in    std_logic
); 
end component;

component FRAME_CHECK 
generic
(
    RX_DATA_WIDTH            : integer := 16;
    USE_COMMA                : integer := 1;
    NONE_MSB_FIRST_DEC       : integer := 0;
    COMMA_DOUBLE_DEC         : integer := 0;
    CHANBOND_SEQ_LEN         : integer := 1;
    WORDS_IN_BRAM            : integer := 256;
    CONFIG_INDEPENDENT_LANES : integer := 0;
    START_OF_PACKET_CHAR     : std_logic_vector := x"55fb";
    COMMA_DOUBLE_CHAR        : std_logic_vector := x"f628";
    MEM_00       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_01       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_02       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_03       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_04       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_05       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_06       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_07       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_08       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_09       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_10       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_11       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_12       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_13       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_14       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_15       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_16       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_17       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_18       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_19       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_20       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_21       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_22       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_23       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_24       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_25       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_26       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_27       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_28       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_29       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_30       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_31       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_32       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_33       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_34       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_35       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_36       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_37       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_38       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_39       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_00      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_01      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_02      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_03      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_04      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_05      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_06      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_07      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000"
);
port
(
    -- User Interface
    RX_DATA                  : in  std_logic_vector((RX_DATA_WIDTH-1) downto 0); 
    RX_ENMCOMMA_ALIGN        : out std_logic;
    RX_ENPCOMMA_ALIGN        : out std_logic;
    RX_ENCHAN_SYNC           : out std_logic; 
    RX_CHANBOND_SEQ          : in  std_logic; 

    -- Control Interface
    INC_IN                   : in std_logic; 
    INC_OUT                  : out std_logic; 
    PATTERN_MATCH_N          : out std_logic;
    RESET_ON_ERROR           : in std_logic; 
    
    -- Error Monitoring
    ERROR_COUNT              : out std_logic_vector(7 downto 0);
    
    -- Track Data
    TRACK_DATA               : out std_logic;

    -- System Interface
    USER_CLK                 : in std_logic;
    SYSTEM_RESET             : in std_logic
  
);
end component;

component MGT_USRCLK_SOURCE_MMCM
generic
(
    MULT                 : real             := 2.0;
    DIVIDE               : integer          := 2;    
    CLK_PERIOD           : real             := 6.4;    
    OUT0_DIVIDE          : real             := 2.0;
    OUT1_DIVIDE          : integer          := 2;
    OUT2_DIVIDE          : integer          := 2;
    OUT3_DIVIDE          : integer          := 2
);
port
( 
    CLK0_OUT                : out std_logic;
    CLK1_OUT                : out std_logic;
    CLK2_OUT                : out std_logic;
    CLK3_OUT                : out std_logic;
    CLK_IN                  : in  std_logic;
    MMCM_LOCKED_OUT         : out std_logic;
    MMCM_RESET_IN           : in  std_logic
);
end component;

component TX_SYNC 
generic
(
    -- Simulation attributes
    SIM_TXPMASETPHASE_SPEEDUP    : integer   := 0 -- Set to 1 to speed up sim reset
);
port
(
    TXENPMAPHASEALIGN       : out std_logic;
    TXPMASETPHASE           : out std_logic;
    TXDLYALIGNDISABLE       : out std_logic;
    TXDLYALIGNRESET         : out std_logic;
    SYNC_DONE               : out std_logic;
    USER_CLK                : in  std_logic;
    RESET                   : in  std_logic
);
end component;


-- Chipscope modules
attribute syn_black_box                : boolean;
attribute syn_noprune                  : boolean;


component data_vio
port
(
    control                 : inout std_logic_vector(35 downto 0);
    clk                     : in    std_logic;
    async_in                : in    std_logic_vector(31 downto 0);
    async_out               : out   std_logic_vector(31 downto 0);
    sync_in                 : in    std_logic_vector(31 downto 0);
    sync_out                : out   std_logic_vector(31 downto 0)
);
end component;
attribute syn_black_box of data_vio : component is TRUE;
attribute syn_noprune of data_vio   : component is TRUE;


component icon
port
(
    control0                : inout std_logic_vector(35 downto 0);
    control1                : inout std_logic_vector(35 downto 0);
    control2                : inout std_logic_vector(35 downto 0);
    control3                : inout std_logic_vector(35 downto 0)
);
end component;
attribute syn_black_box of icon : component is TRUE;
attribute syn_noprune of icon   : component is TRUE;


component ila
port
(
    control                 : inout std_logic_vector(35 downto 0);
    clk                     : in    std_logic;
    trig0                   : in    std_logic_vector(84 downto 0)
);
end component;


attribute syn_black_box of ila : component is TRUE;
attribute syn_noprune of ila   : component is TRUE;


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;
 
    constant ALIGNER_LOOK_INIT : std_logic_vector := "00011111"; 
    constant ALIGNER_LOOK_INCR : std_logic_vector := "00000100";
    constant ALIGNER_LOCK_INCR : std_logic_vector := "010";
    constant ALIGNER_WAIT      : std_logic_vector := "00100000";

    attribute max_fanout : string; 

--************************** Register Declarations ****************************

    signal   gtx0_txresetdone_r              : std_logic;
    signal   gtx0_txresetdone_r2             : std_logic;


--**************************** Wire Declarations ******************************
    -------------------------- MGT Wrapper Wires ------------------------------
    --________________________________________________________________________
    --________________________________________________________________________
    --GTX0   (X0Y2)

    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    signal  gtx0_txcharisk_i                : std_logic_vector(3 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gtx0_txdata_i                   : std_logic_vector(31 downto 0);
    signal  gtx0_txoutclk_i                 : std_logic;
    -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    signal  gtx0_txdlyaligndisable_i        : std_logic;
    signal  gtx0_txdlyalignmonenb_i         : std_logic;
    signal  gtx0_txdlyalignmonitor_i        : std_logic_vector(7 downto 0);
    signal  gtx0_txdlyalignreset_i          : std_logic;
    signal  gtx0_txenpmaphasealign_i        : std_logic;
    signal  gtx0_txpmasetphase_i            : std_logic;
    ----------------------- Transmit Ports - TX PLL Ports ----------------------
    signal  gtx0_gtxtxreset_i               : std_logic;
    signal  gtx0_plltxreset_i               : std_logic;
    signal  gtx0_txplllkdet_i               : std_logic;
    signal  gtx0_txresetdone_i              : std_logic;




    signal  gtx0_tx_system_reset_c          : std_logic;
    signal  gtx0_rx_system_reset_c          : std_logic;
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_ground_vec_i            : std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   : std_logic;
    signal  tied_to_vcc_vec_i               : std_logic_vector(7 downto 0);
    signal  drp_clk_in_i                    : std_logic;
 

    ----------------------------- User Clocks ---------------------------------

    signal  gtx0_txusrclk_i                 : std_logic;
    signal  gtx0_txusrclk2_i                : std_logic;
    signal  txoutclk_mmcm0_locked_i         : std_logic;
    signal  txoutclk_mmcm0_reset_i          : std_logic;
    signal  gtx0_txoutclk_to_mmcm_i         : std_logic;


    ----------------------------- Reference Clocks ----------------------------
    
    signal    q1_clk1_refclk_i                : std_logic;
    signal    q1_clk1_refclk_i_bufg           : std_logic;

    ----------------------- Frame check/gen Module Signals --------------------
    
    signal    gtx0_matchn_i                   : std_logic;
    
    signal    gtx0_txdata_float_i             : std_logic_vector(7 downto 0);
    
    signal    gtx0_track_data_i               : std_logic;
    signal    gtx0_block_sync_i               : std_logic;
    signal    gtx0_error_count_i              : std_logic_vector(7 downto 0);
    signal    gtx0_frame_check_reset_i        : std_logic;
    signal    gtx0_inc_in_i                   : std_logic;
    signal    gtx0_inc_out_i                  : std_logic;
    signal    gtx0_unscrambled_data_i         : std_logic_vector(15 downto 0);

    signal    reset_on_data_error_i           : std_logic;
    signal    track_data_out_i                : std_logic;
 
    
    ------------------------- Sync Module Signals -----------------------------


    signal    gtx0_tx_sync_done_i             : std_logic;
    signal    gtx0_reset_txsync_c             : std_logic;

    ----------------------- Chipscope Signals ---------------------------------

    signal  tx_data_vio_control_i           : std_logic_vector(35 downto 0);
    signal  rx_data_vio_control_i           : std_logic_vector(35 downto 0);
    signal  shared_vio_control_i            : std_logic_vector(35 downto 0);
    signal  ila_control_i                   : std_logic_vector(35 downto 0);
    signal  tx_data_vio_async_in_i          : std_logic_vector(31 downto 0);
    signal  tx_data_vio_sync_in_i           : std_logic_vector(31 downto 0);
    signal  tx_data_vio_async_out_i         : std_logic_vector(31 downto 0);
    signal  tx_data_vio_sync_out_i          : std_logic_vector(31 downto 0);
    signal  rx_data_vio_async_in_i          : std_logic_vector(31 downto 0);
    signal  rx_data_vio_sync_in_i           : std_logic_vector(31 downto 0);
    signal  rx_data_vio_async_out_i         : std_logic_vector(31 downto 0);
    signal  rx_data_vio_sync_out_i          : std_logic_vector(31 downto 0);
    signal  shared_vio_in_i                 : std_logic_vector(31 downto 0);
    signal  shared_vio_out_i                : std_logic_vector(31 downto 0);
    signal  ila_in_i                        : std_logic_vector(84 downto 0);

    signal  gtx0_tx_data_vio_async_in_i     : std_logic_vector(31 downto 0);
    signal  gtx0_tx_data_vio_sync_in_i      : std_logic_vector(31 downto 0);
    signal  gtx0_tx_data_vio_async_out_i    : std_logic_vector(31 downto 0);
    signal  gtx0_tx_data_vio_sync_out_i     : std_logic_vector(31 downto 0);
    signal  gtx0_rx_data_vio_async_in_i     : std_logic_vector(31 downto 0);
    signal  gtx0_rx_data_vio_sync_in_i      : std_logic_vector(31 downto 0);
    signal  gtx0_rx_data_vio_async_out_i    : std_logic_vector(31 downto 0);
    signal  gtx0_rx_data_vio_sync_out_i     : std_logic_vector(31 downto 0);
    signal  gtx0_ila_in_i                   : std_logic_vector(84 downto 0);


    signal    gtxtxreset_i                    : std_logic;
    signal    gtxrxreset_i                    : std_logic;

    signal    user_tx_reset_i                 : std_logic;
    signal    user_rx_reset_i                 : std_logic;
    signal    tx_vio_clk_i                    : std_logic;
    signal    tx_vio_clk_mux_out_i            : std_logic;
    signal    rx_vio_ila_clk_i                : std_logic;
    signal    rx_vio_ila_clk_mux_out_i        : std_logic;

    
--**************************** Main Body of Code *******************************
begin

    --  Static signal Assigments
    tied_to_ground_i                             <= '0';
    tied_to_ground_vec_i                         <= x"0000000000000000";
    tied_to_vcc_i                                <= '1';
    tied_to_vcc_vec_i                            <= x"ff";



    
  

    -----------------------Dedicated GTX Reference Clock Inputs ---------------
    -- The dedicated reference clock inputs you selected in the GUI are implemented using
    -- IBUFDS_GTXE1 instances.
    --
    -- In the UCF file for this example design, you will see that each of
    -- these IBUFDS_GTXE1 instances has been LOCed to a particular set of pins. By LOCing to these
    -- locations, we tell the tools to use the dedicated input buffers to the GTX reference
    -- clock network, rather than general purpose IOs. To select other pins, consult the 
    -- Implementation chapter of UG___, or rerun the wizard.
    --
    -- This network is the highest performace (lowest jitter) option for providing clocks
    -- to the GTX transceivers.
    
    q1_clk1_refclk_ibufds_i : IBUFDS_GTXE1
    port map
    (
        O                               =>      q1_clk1_refclk_i,
        ODIV2                           =>      open,
        CEB                             =>      tied_to_ground_i,
        I                               =>      Q1_CLK1_MGTREFCLK_PAD_P_IN,
        IB                              =>      Q1_CLK1_MGTREFCLK_PAD_N_IN
    );

 

   q1_clk1_refclk_bufg_i : BUFG
    port map
    (
        I                               =>      q1_clk1_refclk_i,
        O                               =>      q1_clk1_refclk_i_bufg
    );



    ----------------------------------- User Clocks ---------------------------
    
    -- The clock resources in this section were added based on userclk source selections on
    -- the Latency, Buffering, and Clocking page of the GUI. A few notes about user clocks:
    -- * The userclk and userclk2 for each GTX datapath (TX and RX) must be phase aligned to 
    --   avoid data errors in the fabric interface whenever the datapath is wider than 10 bits
    -- * To minimize clock resources, you can share clocks between GTXs. GTXs using the same frequency
    --   or multiples of the same frequency can be accomadated using MMCMs. Use caution when
    --   using RXRECCLK as a clock source, however - these clocks can typically only be shared if all
    --   the channels using the clock are receiving data from TX channels that share a reference clock 
    --   source with each other.

    txoutclk_mmcm0_reset_i                       <= not gtx0_txplllkdet_i;
    txoutclk_mmcm0_i : MGT_USRCLK_SOURCE_MMCM
    generic map
    (
        MULT                            =>      8.0,
        DIVIDE                          =>      1,
        CLK_PERIOD                      =>      12.5,
        OUT0_DIVIDE                     =>      8.0,
        OUT1_DIVIDE                     =>      4,
        OUT2_DIVIDE                     =>      1,
        OUT3_DIVIDE                     =>      1
    )
    port map
    (
        CLK0_OUT                        =>      gtx0_txusrclk2_i,
        CLK1_OUT                        =>      gtx0_txusrclk_i,
        CLK2_OUT                        =>      open,
        CLK3_OUT                        =>      open,
        CLK_IN                          =>      gtx0_txoutclk_i,
        MMCM_LOCKED_OUT                 =>      txoutclk_mmcm0_locked_i,
        MMCM_RESET_IN                   =>      txoutclk_mmcm0_reset_i
    );




    ----------------------------- The GTX Wrapper -----------------------------
    
    -- Use the instantiation template in the example directory to add the GTX wrapper to your design.
    -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    -- checker. The GTXs will reset, then attempt to align and transmit data. If channel bonding is 
    -- enabled, bonding should occur after alignment.



    trg_tx_buf_bypass_i : TRG_TX_BUF_BYPASS
    generic map
    (
        WRAPPER_SIM_GTXRESET_SPEEDUP    =>      EXAMPLE_SIM_GTXRESET_SPEEDUP
    )
    port map
    (
  
 
 

        --_____________________________________________________________________
        --_____________________________________________________________________
        --GTX0  (X0Y2)
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        GTX0_RXN_IN                     =>      RXN_IN,
        GTX0_RXP_IN                     =>      RXP_IN,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        GTX0_TXCHARISK_IN               =>      gtx0_txcharisk_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        GTX0_TXDATA_IN                  =>      gtx0_txdata_i,
        GTX0_TXOUTCLK_OUT               =>      gtx0_txoutclk_i,
        GTX0_TXUSRCLK_IN                =>      gtx0_txusrclk_i,
        GTX0_TXUSRCLK2_IN               =>      gtx0_txusrclk2_i,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GTX0_TXN_OUT                    =>      TXN_OUT,
        GTX0_TXP_OUT                    =>      TXP_OUT,
        -------- Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        GTX0_TXDLYALIGNDISABLE_IN       =>      gtx0_txdlyaligndisable_i,
        GTX0_TXDLYALIGNMONENB_IN        =>      gtx0_txdlyalignmonenb_i,
        GTX0_TXDLYALIGNMONITOR_OUT      =>      gtx0_txdlyalignmonitor_i,
        GTX0_TXDLYALIGNRESET_IN         =>      gtx0_txdlyalignreset_i,
        GTX0_TXENPMAPHASEALIGN_IN       =>      gtx0_txenpmaphasealign_i,
        GTX0_TXPMASETPHASE_IN           =>      gtx0_txpmasetphase_i,
        ----------------------- Transmit Ports - TX PLL Ports ----------------------
        GTX0_GTXTXRESET_IN              =>      gtx0_gtxtxreset_i,
        GTX0_MGTREFCLKTX_IN             =>      q1_clk1_refclk_i,
        GTX0_PLLTXRESET_IN              =>      gtx0_plltxreset_i,
        GTX0_TXPLLLKDET_OUT             =>      gtx0_txplllkdet_i,
        GTX0_TXRESETDONE_OUT            =>      gtx0_txresetdone_i


    );


    ------------------------------ TXSYNC module ------------------------------
    -- The TXSYNC module performs phase synchronization for all the active TX datapaths. It
    -- waits for the user clocks to be stable, then drives the phase align signals on each
    -- GTX. When phase synchronization is complete, it asserts SYNC_DONE
    
    -- Include the TX_SYNC module in your own design to perform phase synchronization if
    -- your protocol bypasses the TX Buffers

  
    
    gtx0_reset_txsync_c  <=  not gtx0_txresetdone_r2;  

    -- SIM_TXPMASETPHASE_SPEEDUP is a simulation only attribute and MUST be set to 0 
    -- during implementation      
    gtx0_txsync_i : TX_SYNC
    generic map
    (
        SIM_TXPMASETPHASE_SPEEDUP       =>      EXAMPLE_SIM_GTXRESET_SPEEDUP
    )
    port map
    (
        TXENPMAPHASEALIGN               =>      gtx0_txenpmaphasealign_i,
        TXPMASETPHASE                   =>      gtx0_txpmasetphase_i,
        TXDLYALIGNDISABLE               =>      gtx0_txdlyaligndisable_i,
        TXDLYALIGNRESET                 =>      gtx0_txdlyalignreset_i,
        SYNC_DONE                       =>      gtx0_tx_sync_done_i,
        USER_CLK                        =>      gtx0_txusrclk2_i,
        RESET                           =>      gtx0_reset_txsync_c
    );



    -------------------------- User Module Resets -----------------------------
    -- All the User Modules i.e. FRAME_GEN, FRAME_CHECK and the sync modules
    -- are held in reset till the RESETDONE goes high. 
    -- The RESETDONE is registered a couple of times on USRCLK2 and connected 
    -- to the reset of the modules
    
    process( gtx0_txusrclk2_i,gtx0_txresetdone_i)
    begin
        if(gtx0_txresetdone_i = '0') then
            gtx0_txresetdone_r  <= '0'   after DLY;
            gtx0_txresetdone_r2 <= '0'   after DLY;
        elsif(gtx0_txusrclk2_i'event and gtx0_txusrclk2_i = '1') then
            gtx0_txresetdone_r  <= gtx0_txresetdone_i   after DLY;
            gtx0_txresetdone_r2 <= gtx0_txresetdone_r   after DLY;
        end if;
    end process;


    ------------------------------ Frame Generators ---------------------------
    -- The example design uses Block RAM based frame generators to provide test
    -- data to the GTXs for transmission. By default the frame generators are 
    -- loaded with an incrementing data sequence that includes commas/alignment
    -- characters for alignment. If your protocol uses channel bonding, the 
    -- frame generator will also be preloaded with a channel bonding sequence.
    
    -- You can modify the data transmitted by changing the INIT values of the frame
    -- generator in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.

    gtx0_frame_gen : FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        MEM_00                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_01                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_02                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_03                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_04                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_05                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_06                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_07                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_08                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_09                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_0A                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_0B                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_0C                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_0D                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_0E                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_0F                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_10                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_11                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_12                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_13                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_14                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_15                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_16                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_17                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_18                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_19                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_1A                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_1B                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_1C                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_1D                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_1E                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_1F                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_20                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_21                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_22                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_23                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_24                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_25                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_26                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_27                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_28                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_29                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_2A                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_2B                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_2C                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_2D                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_2E                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_2F                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_30                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_31                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_32                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_33                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_34                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_35                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_36                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_37                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_38                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_39                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_3A                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_3B                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEM_3C                  =>  x"1e1d1c1b1a191817161514131211100f0e0d0c0b0a0908bc0706050403020100",
        MEM_3D                  =>  x"3e3d3c3b3a393837363534333231302f2e2d2c2b2a292827262524232221201f",
        MEM_3E                  =>  x"5e5d5c5b5a595857565554535251504f4e4d4c4b4a494847464544434241403f",
        MEM_3F                  =>  x"7e7d7c7b7a797877767574737271706f6e6d6c6b6a696867666564636261605f",
        MEMP_00                  =>  x"0000000000000000000000000000010000000000000000000000000000000100",
        MEMP_01                  =>  x"0000000000000000000000000000010000000000000000000000000000000100",
        MEMP_02                  =>  x"0000000000000000000000000000010000000000000000000000000000000100",
        MEMP_03                  =>  x"0000000000000000000000000000010000000000000000000000000000000100",
        MEMP_04                  =>  x"0000000000000000000000000000010000000000000000000000000000000100",
        MEMP_05                  =>  x"0000000000000000000000000000010000000000000000000000000000000100",
        MEMP_06                  =>  x"0000000000000000000000000000010000000000000000000000000000000100",
        MEMP_07                  =>  x"0000000000000000000000000000010000000000000000000000000000000100"
    )
    port map
    (
        -- User Interface
        TX_DATA(39 downto 32)           =>      gtx0_txdata_float_i,
        TX_DATA(31 downto 0)            =>      gtx0_txdata_i,
        TX_CHARISK(3 downto 0)          =>      gtx0_txcharisk_i,
        -- System Interface
        USER_CLK                        =>      gtx0_txusrclk2_i,
        SYSTEM_RESET                    =>      gtx0_tx_system_reset_c
    );
    


    ---------------------------------- Frame Checkers -------------------------
    -- The example design uses Block RAM based frame checkers to verify incoming  
    -- data. By default the frame generators are loaded with a data sequence that 
    -- matches the outgoing sequence of the frame generators for the TX ports.
    
    -- You can modify the expected data sequence by changing the INIT values of the frame
    -- checkers in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.
    
    -- When the frame checker receives data, it attempts to synchronise to the 
    -- incoming pattern by looking for the first sequence in the pattern. Once it 
    -- finds the first sequence, it increments through the sequence, and indicates an 
    -- error whenever the next value received does not match the expected value.

     -- This GTX is not active.The match port for pattern checker of this GTX is tied off
    gtx0_matchn_i                                <= '0';





    ----------------------------- Chipscope Connections -----------------------
    -- When the example design is run in hardware, it uses chipscope to allow the
    -- example design and GTX wrapper to be controlled and monitored. The 
    -- EXAMPLE_USE_CHIPSCOPE parameter allows chipscope to be removed for simulation.
    
chipscope : if EXAMPLE_USE_CHIPSCOPE = 1 generate
    
    
    -- Shared VIO for all transievers 
    shared_vio_i : data_vio
    port map
    (
        control                         =>      shared_vio_control_i,
        clk                             =>      tied_to_ground_i,
        async_in                        =>      shared_vio_in_i,
        async_out                       =>      shared_vio_out_i,
        sync_in                         =>      tied_to_ground_vec_i(31 downto 0),
        sync_out                        =>      open
    );
    
    -- ICON for all VIOs 
    i_icon : icon
    port map
    (
        control0                        =>      shared_vio_control_i,
        control1                        =>      tx_data_vio_control_i,
        control2                        =>      rx_data_vio_control_i,
        control3                        =>      ila_control_i
    );

    
    -- TX VIO 
    tx_data_vio_i : data_vio
    port map
    (
        control                         =>      tx_data_vio_control_i,
        clk                             =>      gtx0_txusrclk2_i,
        async_in                        =>      tx_data_vio_async_in_i,
        async_out                       =>      tx_data_vio_async_out_i,
        sync_in                         =>      tx_data_vio_sync_in_i,
        sync_out                        =>      tx_data_vio_sync_out_i
    );
    
    -- RX VIO 
    rx_data_vio_i : data_vio
    port map
    (
        control                         =>      rx_data_vio_control_i,
        clk                             =>      gtx0_txusrclk2_i,
        async_in                        =>      rx_data_vio_async_in_i,
        async_out                       =>      rx_data_vio_async_out_i,
        sync_in                         =>      rx_data_vio_sync_in_i,
        sync_out                        =>      rx_data_vio_sync_out_i
    );
    
    -- RX ILA
    ila_i : ila
    port map
    (
        control                         =>      ila_control_i,
        clk                             =>      gtx0_txusrclk2_i,
        trig0                           =>      ila_in_i
    );



    -- assign resets for frame_gen modules
    gtx0_tx_system_reset_c                       <= not gtx0_tx_sync_done_i or user_tx_reset_i;
    -- assign resets for frame_check modules

    gtx0_gtxtxreset_i                            <= gtxtxreset_i;

    -- Shared VIO Outputs
    gtxtxreset_i                                 <= shared_vio_out_i(31);
    user_tx_reset_i                              <= shared_vio_out_i(30);
    user_rx_reset_i                              <= shared_vio_out_i(29);

    -- Shared VIO Inputs
    shared_vio_in_i(31 downto 0)                 <= "00000000000000000000000000000000";

    -- Chipscope connections on GTX 0
    gtx0_tx_data_vio_async_in_i(31)              <= gtx0_txplllkdet_i;
    gtx0_tx_data_vio_async_in_i(30)              <= gtx0_txresetdone_i;
    gtx0_tx_data_vio_async_in_i(29 downto 22)    <= gtx0_txdlyalignmonitor_i;
    gtx0_tx_data_vio_async_in_i(21 downto 0)     <= "0000000000000000000000";
    gtx0_tx_data_vio_sync_in_i(31 downto 0)      <= "00000000000000000000000000000000";
    gtx0_plltxreset_i                            <= tx_data_vio_async_out_i(31);
    gtx0_txdlyalignmonenb_i                      <= tx_data_vio_async_out_i(30);
    gtx0_rx_data_vio_async_in_i(31 downto 0)     <= "00000000000000000000000000000000";
    gtx0_rx_data_vio_sync_in_i(31 downto 0)      <= "00000000000000000000000000000000";
    gtx0_ila_in_i(84 downto 77)                  <= gtx0_error_count_i;
    gtx0_ila_in_i(76 downto 0)                   <= "00000000000000000000000000000000000000000000000000000000000000000000000000000";



    tx_data_vio_async_in_i              <=      gtx0_tx_data_vio_async_in_i;


    tx_data_vio_sync_in_i               <=      gtx0_tx_data_vio_sync_in_i;

    rx_data_vio_async_in_i              <=      gtx0_rx_data_vio_async_in_i;


    rx_data_vio_sync_in_i               <=      gtx0_rx_data_vio_sync_in_i;


    ila_in_i                            <=      gtx0_ila_in_i;


end generate chipscope;


no_chipscope : if EXAMPLE_USE_CHIPSCOPE = 0 generate

    -- If Chipscope is not being used, drive GTX reset signal
    -- from the top level ports
    gtx0_gtxtxreset_i                            <= GTXTXRESET_IN;

    -- assign resets for frame_gen modules
    gtx0_tx_system_reset_c                       <= not gtx0_tx_sync_done_i;
    -- assign resets for frame_check modules

    gtxtxreset_i                                 <= tied_to_ground_i;
    user_tx_reset_i                              <= tied_to_ground_i;
    user_rx_reset_i                              <= tied_to_ground_i;
    gtx0_plltxreset_i                            <= tied_to_ground_i;
    gtx0_txdlyalignmonenb_i                      <= tied_to_ground_i;



end generate no_chipscope;


end RTL;


