///////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 1.8
//  \   \         Application : Virtex-6 FPGA GTX Transceiver Wizard
//  /   /         Filename : snap12_t20r20.v
// /___/   /\     
// \   \  /  \ 
//  \___\/\___\
//
//
// Module SNAP12_T20R20 (a GTX Wrapper)
// Generated by Xilinx Virtex-6 FPGA GTX Transceiver Wizard
// 

`timescale 1ns / 1ps


//***************************** Entity Declaration ****************************

(* CORE_GENERATION_INFO = "SNAP12_T20R20,v6_gtxwizard_v1_8,{protocol_file=aurora_2byte_single_lane}" *)
module SNAP12_T20R20 #
(
    // Simulation attributes
    parameter   WRAPPER_SIM_GTXRESET_SPEEDUP    = 0    // Set to 1 to speed up sim reset
)
(
    input gtx_wait,
    output [11:0] rxdv_snapr, rxcomma_snapr, // my RxDV and Comma
    output [11:0] check_ok_snapr, check_bad_snapr, good_byte, bad_byte, lost_byte,
    output [31:0] errcount0,
    output [31:0] errcount1,
    output [31:0] errcount2,
    output [31:0] errcount3,
    output [31:0] errcount4,
    output [31:0] errcount5,
    output [31:0] errcount6,
    output [31:0] errcount7,
    output [31:0] errcount8,
    output [31:0] errcount9,
    output [31:0] errcount10,
    output [31:0] errcount11,
    output [15:0] GTXi_RXDATA_OUT,  // select just ONE gtx data to monitor...
    output  [1:0] GTXi_RXK_OUT,     // select the K that goes with it

    //_________________________________________________________________________
    //_________________________________________________________________________
    //GTX0  (X0Y0)
    //---------------------- Loopback and Powerdown Ports ----------------------
//jg    input   [1:0]   GTX0_RXPOWERDOWN_IN,
//jg    input   [1:0]   GTX0_TXPOWERDOWN_IN,
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg    output  [1:0]   GTX0_RXCHARISCOMMA_OUT,
//jg    output  [1:0]   GTX0_RXDISPERR_OUT,
//jg    output  [1:0]   GTX0_RXNOTINTABLE_OUT,
    //----------------- Receive Ports - Clock Correction Ports -----------------
    output  [2:0]   GTX0_RXCLKCORCNT_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          GTX0_RXBYTEREALIGN_OUT,
    output          GTX0_RXCOMMADET_OUT,      //jg: useful?
    input           GTX0_RXENMCOMMAALIGN_IN,
    input           GTX0_RXENPCOMMAALIGN_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
//jg    output  [15:0]  GTX0_RXDATA_OUT,
    input           GTX0_RXRESET_IN,
    input           GTX0_RXUSRCLK2_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input           GTX0_RXCDRRESET_IN,
    input           GTX0_RXN_IN,
    input           GTX0_RXP_IN,
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg    output  [2:0]   GTX0_RXBUFSTATUS_OUT,
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    output  [1:0]   GTX0_RXLOSSOFSYNC_OUT,
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    input           GTX0_GTXRXRESET_IN,
    input           GTX0_MGTREFCLKRX_IN,
    input           GTX0_PLLRXRESET_IN,
    output          GTX0_RXPLLLKDET_OUT,
    output          GTX0_RXRESETDONE_OUT,
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    output          GTX0_RXVALID_OUT,         //jg: useful?
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           GTX0_RXPOLARITY_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [64:0]  GTX0_SEED_IN,
    input   [64:0]  GTX0_RXSEED,
    output          GTX0_TXOUTCLK_OUT,
    input           GTX0_TXRESET_IN,
    input           GTX0_TXUSRCLK2_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GTX0_TXN_OUT,
    output          GTX0_TXP_OUT,
    input           gtx0_force_error,
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    input           GTX0_TXDLYALIGNDISABLE_IN,
    input           GTX0_TXDLYALIGNMONENB_IN,
    output  [7:0]   GTX0_TXDLYALIGNMONITOR_OUT,
    input           GTX0_TXDLYALIGNRESET_IN,
    input           GTX0_TXENPMAPHASEALIGN_IN,
    input           GTX0_TXPMASETPHASE_IN,
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    input           GTX0_GTXTXRESET_IN,
    output          GTX0_TXRESETDONE_OUT,

    //_________________________________________________________________________
    //_________________________________________________________________________
    //GTX1  (X0Y1)
    //---------------------- Loopback and Powerdown Ports ----------------------
//jg    input   [1:0]   GTX1_RXPOWERDOWN_IN,
//jg    input   [1:0]   GTX1_TXPOWERDOWN_IN,
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg    output  [1:0]   GTX1_RXCHARISCOMMA_OUT,
//jg    output  [1:0]   GTX1_RXDISPERR_OUT,
//jg    output  [1:0]   GTX1_RXNOTINTABLE_OUT,
    //----------------- Receive Ports - Clock Correction Ports -----------------
    output  [2:0]   GTX1_RXCLKCORCNT_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          GTX1_RXBYTEREALIGN_OUT,
    output          GTX1_RXCOMMADET_OUT,
    input           GTX1_RXENMCOMMAALIGN_IN,
    input           GTX1_RXENPCOMMAALIGN_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
//jg    output  [15:0]  GTX1_RXDATA_OUT,
    input           GTX1_RXRESET_IN,
    input           GTX1_RXUSRCLK2_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input           GTX1_RXCDRRESET_IN,
    input           GTX1_RXN_IN,
    input           GTX1_RXP_IN,
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg    output  [2:0]   GTX1_RXBUFSTATUS_OUT,
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    output  [1:0]   GTX1_RXLOSSOFSYNC_OUT,
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    input           GTX1_GTXRXRESET_IN,
    input           GTX1_MGTREFCLKRX_IN,
    input           GTX1_PLLRXRESET_IN,
    output          GTX1_RXPLLLKDET_OUT,
    output          GTX1_RXRESETDONE_OUT,
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    output          GTX1_RXVALID_OUT,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           GTX1_RXPOLARITY_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [64:0]  GTX1_SEED_IN,
    input   [64:0]  GTX1_RXSEED,
    output          GTX1_TXOUTCLK_OUT,
    input           GTX1_TXRESET_IN,
    input           GTX1_TXUSRCLK2_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GTX1_TXN_OUT,
    output          GTX1_TXP_OUT,
    input           gtx1_force_error,
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    input           GTX1_TXDLYALIGNDISABLE_IN,
    input           GTX1_TXDLYALIGNMONENB_IN,
    output  [7:0]   GTX1_TXDLYALIGNMONITOR_OUT,
    input           GTX1_TXDLYALIGNRESET_IN,
    input           GTX1_TXENPMAPHASEALIGN_IN,
    input           GTX1_TXPMASETPHASE_IN,
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    input           GTX1_GTXTXRESET_IN,
    output          GTX1_TXRESETDONE_OUT,

    //_________________________________________________________________________
    //_________________________________________________________________________
    //GTX2  (X0Y2)
    //---------------------- Loopback and Powerdown Ports ----------------------
//jg    input   [1:0]   GTX2_RXPOWERDOWN_IN,
//jg    input   [1:0]   GTX2_TXPOWERDOWN_IN,
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg    output  [1:0]   GTX2_RXCHARISCOMMA_OUT,
//jg    output  [1:0]   GTX2_RXDISPERR_OUT,
//jg    output  [1:0]   GTX2_RXNOTINTABLE_OUT,
    //----------------- Receive Ports - Clock Correction Ports -----------------
    output  [2:0]   GTX2_RXCLKCORCNT_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          GTX2_RXBYTEREALIGN_OUT,
    output          GTX2_RXCOMMADET_OUT,
    input           GTX2_RXENMCOMMAALIGN_IN,
    input           GTX2_RXENPCOMMAALIGN_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
//jg    output  [15:0]  GTX2_RXDATA_OUT,
    input           GTX2_RXRESET_IN,
    input           GTX2_RXUSRCLK2_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input           GTX2_RXCDRRESET_IN,
    input           GTX2_RXN_IN,
    input           GTX2_RXP_IN,
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg    output  [2:0]   GTX2_RXBUFSTATUS_OUT,
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    output  [1:0]   GTX2_RXLOSSOFSYNC_OUT,
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    input           GTX2_GTXRXRESET_IN,
    input           GTX2_MGTREFCLKRX_IN,
    input           GTX2_PLLRXRESET_IN,
    output          GTX2_RXPLLLKDET_OUT,
    output          GTX2_RXRESETDONE_OUT,
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    output          GTX2_RXVALID_OUT,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           GTX2_RXPOLARITY_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [64:0]  GTX2_SEED_IN,
    input   [64:0]  GTX2_RXSEED,
    output          GTX2_TXOUTCLK_OUT,
    input           GTX2_TXRESET_IN,
    input           GTX2_TXUSRCLK2_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GTX2_TXN_OUT,
    output          GTX2_TXP_OUT,
    input           gtx2_force_error,
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    input           GTX2_TXDLYALIGNDISABLE_IN,
    input           GTX2_TXDLYALIGNMONENB_IN,
    output  [7:0]   GTX2_TXDLYALIGNMONITOR_OUT,
    input           GTX2_TXDLYALIGNRESET_IN,
    input           GTX2_TXENPMAPHASEALIGN_IN,
    input           GTX2_TXPMASETPHASE_IN,
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    input           GTX2_GTXTXRESET_IN,
    output          GTX2_TXRESETDONE_OUT,

    //_________________________________________________________________________
    //_________________________________________________________________________
    //GTX3  (X0Y3)
    //---------------------- Loopback and Powerdown Ports ----------------------
//jg    input   [1:0]   GTX3_RXPOWERDOWN_IN,
//jg    input   [1:0]   GTX3_TXPOWERDOWN_IN,
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg    output  [1:0]   GTX3_RXCHARISCOMMA_OUT,
//jg    output  [1:0]   GTX3_RXDISPERR_OUT,
//jg    output  [1:0]   GTX3_RXNOTINTABLE_OUT,
    //----------------- Receive Ports - Clock Correction Ports -----------------
    output  [2:0]   GTX3_RXCLKCORCNT_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          GTX3_RXBYTEREALIGN_OUT,
    output          GTX3_RXCOMMADET_OUT,
    input           GTX3_RXENMCOMMAALIGN_IN,
    input           GTX3_RXENPCOMMAALIGN_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
//jg    output  [15:0]  GTX3_RXDATA_OUT,
    input           GTX3_RXRESET_IN,
    input           GTX3_RXUSRCLK2_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input           GTX3_RXCDRRESET_IN,
    input           GTX3_RXN_IN,
    input           GTX3_RXP_IN,
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg    output  [2:0]   GTX3_RXBUFSTATUS_OUT,
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    output  [1:0]   GTX3_RXLOSSOFSYNC_OUT,
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    input           GTX3_GTXRXRESET_IN,
    input           GTX3_MGTREFCLKRX_IN,
    input           GTX3_PLLRXRESET_IN,
    output          GTX3_RXPLLLKDET_OUT,
    output          GTX3_RXRESETDONE_OUT,
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    output          GTX3_RXVALID_OUT,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           GTX3_RXPOLARITY_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [64:0]  GTX3_SEED_IN,
    input   [64:0]  GTX3_RXSEED,
    output          GTX3_TXOUTCLK_OUT,
    input           GTX3_TXRESET_IN,
    input           GTX3_TXUSRCLK2_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GTX3_TXN_OUT,
    output          GTX3_TXP_OUT,
    input           gtx3_force_error,
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    input           GTX3_TXDLYALIGNDISABLE_IN,
    input           GTX3_TXDLYALIGNMONENB_IN,
    output  [7:0]   GTX3_TXDLYALIGNMONITOR_OUT,
    input           GTX3_TXDLYALIGNRESET_IN,
    input           GTX3_TXENPMAPHASEALIGN_IN,
    input           GTX3_TXPMASETPHASE_IN,
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    input           GTX3_GTXTXRESET_IN,
    output          GTX3_TXRESETDONE_OUT,

    //_________________________________________________________________________
    //_________________________________________________________________________
    //GTX4  (X0Y4)
    //---------------------- Loopback and Powerdown Ports ----------------------
//jg    input   [1:0]   GTX4_RXPOWERDOWN_IN,
//jg    input   [1:0]   GTX4_TXPOWERDOWN_IN,
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg    output  [1:0]   GTX4_RXCHARISCOMMA_OUT,
//jg    output  [1:0]   GTX4_RXDISPERR_OUT,
//jg    output  [1:0]   GTX4_RXNOTINTABLE_OUT,
    //----------------- Receive Ports - Clock Correction Ports -----------------
    output  [2:0]   GTX4_RXCLKCORCNT_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          GTX4_RXBYTEREALIGN_OUT,
    output          GTX4_RXCOMMADET_OUT,
    input           GTX4_RXENMCOMMAALIGN_IN,
    input           GTX4_RXENPCOMMAALIGN_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
//jg    output  [15:0]  GTX4_RXDATA_OUT,
    input           GTX4_RXRESET_IN,
    input           GTX4_RXUSRCLK2_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input           GTX4_RXCDRRESET_IN,
    input           GTX4_RXN_IN,
    input           GTX4_RXP_IN,
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg    output  [2:0]   GTX4_RXBUFSTATUS_OUT,
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    output  [1:0]   GTX4_RXLOSSOFSYNC_OUT,
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    input           GTX4_GTXRXRESET_IN,
    input           GTX4_MGTREFCLKRX_IN,
    input           GTX4_PLLRXRESET_IN,
    output          GTX4_RXPLLLKDET_OUT,
    output          GTX4_RXRESETDONE_OUT,
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    output          GTX4_RXVALID_OUT,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           GTX4_RXPOLARITY_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [64:0]  GTX4_SEED_IN,
    input   [64:0]  GTX4_RXSEED,
    output          GTX4_TXOUTCLK_OUT,
    input           GTX4_TXRESET_IN,
    input           GTX4_TXUSRCLK2_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GTX4_TXN_OUT,
    output          GTX4_TXP_OUT,
    input           gtx4_force_error,
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    input           GTX4_TXDLYALIGNDISABLE_IN,
    input           GTX4_TXDLYALIGNMONENB_IN,
    output  [7:0]   GTX4_TXDLYALIGNMONITOR_OUT,
    input           GTX4_TXDLYALIGNRESET_IN,
    input           GTX4_TXENPMAPHASEALIGN_IN,
    input           GTX4_TXPMASETPHASE_IN,
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    input           GTX4_GTXTXRESET_IN,
    output          GTX4_TXRESETDONE_OUT,

    //_________________________________________________________________________
    //_________________________________________________________________________
    //GTX5  (X0Y5)
    //---------------------- Loopback and Powerdown Ports ----------------------
//jg    input   [1:0]   GTX5_RXPOWERDOWN_IN,
//jg    input   [1:0]   GTX5_TXPOWERDOWN_IN,
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg    output  [1:0]   GTX5_RXCHARISCOMMA_OUT,
//jg    output  [1:0]   GTX5_RXDISPERR_OUT,
//jg    output  [1:0]   GTX5_RXNOTINTABLE_OUT,
    //----------------- Receive Ports - Clock Correction Ports -----------------
    output  [2:0]   GTX5_RXCLKCORCNT_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          GTX5_RXBYTEREALIGN_OUT,
    output          GTX5_RXCOMMADET_OUT,
    input           GTX5_RXENMCOMMAALIGN_IN,
    input           GTX5_RXENPCOMMAALIGN_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
//jg    output  [15:0]  GTX5_RXDATA_OUT,
    input           GTX5_RXRESET_IN,
    input           GTX5_RXUSRCLK2_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input           GTX5_RXCDRRESET_IN,
    input           GTX5_RXN_IN,
    input           GTX5_RXP_IN,
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg    output  [2:0]   GTX5_RXBUFSTATUS_OUT,
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    output  [1:0]   GTX5_RXLOSSOFSYNC_OUT,
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    input           GTX5_GTXRXRESET_IN,
    input           GTX5_MGTREFCLKRX_IN,
    input           GTX5_PLLRXRESET_IN,
    output          GTX5_RXPLLLKDET_OUT,
    output          GTX5_RXRESETDONE_OUT,
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    output          GTX5_RXVALID_OUT,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           GTX5_RXPOLARITY_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [64:0]  GTX5_SEED_IN,
    input   [64:0]  GTX5_RXSEED,
    output          GTX5_TXOUTCLK_OUT,
    input           GTX5_TXRESET_IN,
    input           GTX5_TXUSRCLK2_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GTX5_TXN_OUT,
    output          GTX5_TXP_OUT,
    input           gtx5_force_error,
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    input           GTX5_TXDLYALIGNDISABLE_IN,
    input           GTX5_TXDLYALIGNMONENB_IN,
    output  [7:0]   GTX5_TXDLYALIGNMONITOR_OUT,
    input           GTX5_TXDLYALIGNRESET_IN,
    input           GTX5_TXENPMAPHASEALIGN_IN,
    input           GTX5_TXPMASETPHASE_IN,
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    input           GTX5_GTXTXRESET_IN,
    output          GTX5_TXRESETDONE_OUT,

    //_________________________________________________________________________
    //_________________________________________________________________________
    //GTX6  (X0Y6)
    //---------------------- Loopback and Powerdown Ports ----------------------
//jg    input   [1:0]   GTX6_RXPOWERDOWN_IN,
//jg    input   [1:0]   GTX6_TXPOWERDOWN_IN,
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg    output  [1:0]   GTX6_RXCHARISCOMMA_OUT,
//jg    output  [1:0]   GTX6_RXDISPERR_OUT,
//jg    output  [1:0]   GTX6_RXNOTINTABLE_OUT,
    //----------------- Receive Ports - Clock Correction Ports -----------------
    output  [2:0]   GTX6_RXCLKCORCNT_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          GTX6_RXBYTEREALIGN_OUT,
    output          GTX6_RXCOMMADET_OUT,
    input           GTX6_RXENMCOMMAALIGN_IN,
    input           GTX6_RXENPCOMMAALIGN_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
//jg    output  [15:0]  GTX6_RXDATA_OUT,
    input           GTX6_RXRESET_IN,
    input           GTX6_RXUSRCLK2_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input           GTX6_RXCDRRESET_IN,
    input           GTX6_RXN_IN,
    input           GTX6_RXP_IN,
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg    output  [2:0]   GTX6_RXBUFSTATUS_OUT,
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    output  [1:0]   GTX6_RXLOSSOFSYNC_OUT,
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    input           GTX6_GTXRXRESET_IN,
    input           GTX6_MGTREFCLKRX_IN,
    input           GTX6_PLLRXRESET_IN,
    output          GTX6_RXPLLLKDET_OUT,
    output          GTX6_RXRESETDONE_OUT,
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    output          GTX6_RXVALID_OUT,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           GTX6_RXPOLARITY_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [64:0]  GTX6_SEED_IN,
    input   [64:0]  GTX6_RXSEED,
    output          GTX6_TXOUTCLK_OUT,
    input           GTX6_TXRESET_IN,
    input           GTX6_TXUSRCLK2_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GTX6_TXN_OUT,
    output          GTX6_TXP_OUT,
    input           gtx6_force_error,
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    input           GTX6_TXDLYALIGNDISABLE_IN,
    input           GTX6_TXDLYALIGNMONENB_IN,
    output  [7:0]   GTX6_TXDLYALIGNMONITOR_OUT,
    input           GTX6_TXDLYALIGNRESET_IN,
    input           GTX6_TXENPMAPHASEALIGN_IN,
    input           GTX6_TXPMASETPHASE_IN,
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    input           GTX6_GTXTXRESET_IN,
    output          GTX6_TXRESETDONE_OUT,

    //_________________________________________________________________________
    //_________________________________________________________________________
    //GTX7  (X0Y7)
    //---------------------- Loopback and Powerdown Ports ----------------------
//jg    input   [1:0]   GTX7_RXPOWERDOWN_IN,
//jg    input   [1:0]   GTX7_TXPOWERDOWN_IN,
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg    output  [1:0]   GTX7_RXCHARISCOMMA_OUT,
//jg    output  [1:0]   GTX7_RXDISPERR_OUT,
//jg    output  [1:0]   GTX7_RXNOTINTABLE_OUT,
    //----------------- Receive Ports - Clock Correction Ports -----------------
    output  [2:0]   GTX7_RXCLKCORCNT_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          GTX7_RXBYTEREALIGN_OUT,
    output          GTX7_RXCOMMADET_OUT,
    input           GTX7_RXENMCOMMAALIGN_IN,
    input           GTX7_RXENPCOMMAALIGN_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
//jg    output  [15:0]  GTX7_RXDATA_OUT,
    input           GTX7_RXRESET_IN,
    input           GTX7_RXUSRCLK2_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input           GTX7_RXCDRRESET_IN,
    input           GTX7_RXN_IN,
    input           GTX7_RXP_IN,
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg    output  [2:0]   GTX7_RXBUFSTATUS_OUT,
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    output  [1:0]   GTX7_RXLOSSOFSYNC_OUT,
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    input           GTX7_GTXRXRESET_IN,
    input           GTX7_MGTREFCLKRX_IN,
    input           GTX7_PLLRXRESET_IN,
    output          GTX7_RXPLLLKDET_OUT,
    output          GTX7_RXRESETDONE_OUT,
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    output          GTX7_RXVALID_OUT,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           GTX7_RXPOLARITY_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [64:0]  GTX7_SEED_IN,
    input   [64:0]  GTX7_RXSEED,
    output          GTX7_TXOUTCLK_OUT,
    input           GTX7_TXRESET_IN,
    input           GTX7_TXUSRCLK2_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GTX7_TXN_OUT,
    output          GTX7_TXP_OUT,
    input           gtx7_force_error,
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    input           GTX7_TXDLYALIGNDISABLE_IN,
    input           GTX7_TXDLYALIGNMONENB_IN,
    output  [7:0]   GTX7_TXDLYALIGNMONITOR_OUT,
    input           GTX7_TXDLYALIGNRESET_IN,
    input           GTX7_TXENPMAPHASEALIGN_IN,
    input           GTX7_TXPMASETPHASE_IN,
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    input           GTX7_GTXTXRESET_IN,
    output          GTX7_TXRESETDONE_OUT,

    //_________________________________________________________________________
    //_________________________________________________________________________
    //GTX8  (X0Y8)
    //---------------------- Loopback and Powerdown Ports ----------------------
//jg    input   [1:0]   GTX8_RXPOWERDOWN_IN,
//jg    input   [1:0]   GTX8_TXPOWERDOWN_IN,
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg    output  [1:0]   GTX8_RXCHARISCOMMA_OUT,
//jg    output  [1:0]   GTX8_RXDISPERR_OUT,
//jg    output  [1:0]   GTX8_RXNOTINTABLE_OUT,
    //----------------- Receive Ports - Clock Correction Ports -----------------
    output  [2:0]   GTX8_RXCLKCORCNT_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          GTX8_RXBYTEREALIGN_OUT,
    output          GTX8_RXCOMMADET_OUT,
    input           GTX8_RXENMCOMMAALIGN_IN,
    input           GTX8_RXENPCOMMAALIGN_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
//jg    output  [15:0]  GTX8_RXDATA_OUT,
    input           GTX8_RXRESET_IN,
    input           GTX8_RXUSRCLK2_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input           GTX8_RXCDRRESET_IN,
    input           GTX8_RXN_IN,
    input           GTX8_RXP_IN,
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg    output  [2:0]   GTX8_RXBUFSTATUS_OUT,
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    output  [1:0]   GTX8_RXLOSSOFSYNC_OUT,
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    input           GTX8_GTXRXRESET_IN,
    input           GTX8_MGTREFCLKRX_IN,
    input           GTX8_PLLRXRESET_IN,
    output          GTX8_RXPLLLKDET_OUT,
    output          GTX8_RXRESETDONE_OUT,
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    output          GTX8_RXVALID_OUT,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           GTX8_RXPOLARITY_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [64:0]  GTX8_SEED_IN,
    input   [64:0]  GTX8_RXSEED,
    output          GTX8_TXOUTCLK_OUT,
    input           GTX8_TXRESET_IN,
    input           GTX8_TXUSRCLK2_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GTX8_TXN_OUT,
    output          GTX8_TXP_OUT,
    input           gtx8_force_error,
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    input           GTX8_TXDLYALIGNDISABLE_IN,
    input           GTX8_TXDLYALIGNMONENB_IN,
    output  [7:0]   GTX8_TXDLYALIGNMONITOR_OUT,
    input           GTX8_TXDLYALIGNRESET_IN,
    input           GTX8_TXENPMAPHASEALIGN_IN,
    input           GTX8_TXPMASETPHASE_IN,
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    input           GTX8_GTXTXRESET_IN,
    output          GTX8_TXRESETDONE_OUT,

    //_________________________________________________________________________
    //_________________________________________________________________________
    //GTX9  (X0Y9)
    //---------------------- Loopback and Powerdown Ports ----------------------
//jg    input   [1:0]   GTX9_RXPOWERDOWN_IN,
//jg    input   [1:0]   GTX9_TXPOWERDOWN_IN,
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg    output  [1:0]   GTX9_RXCHARISCOMMA_OUT,
//jg    output  [1:0]   GTX9_RXDISPERR_OUT,
//jg    output  [1:0]   GTX9_RXNOTINTABLE_OUT,
    //----------------- Receive Ports - Clock Correction Ports -----------------
    output  [2:0]   GTX9_RXCLKCORCNT_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          GTX9_RXBYTEREALIGN_OUT,
    output          GTX9_RXCOMMADET_OUT,
    input           GTX9_RXENMCOMMAALIGN_IN,
    input           GTX9_RXENPCOMMAALIGN_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
//jg    output  [15:0]  GTX9_RXDATA_OUT,
    input           GTX9_RXRESET_IN,
    input           GTX9_RXUSRCLK2_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input           GTX9_RXCDRRESET_IN,
    input           GTX9_RXN_IN,
    input           GTX9_RXP_IN,
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg    output  [2:0]   GTX9_RXBUFSTATUS_OUT,
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    output  [1:0]   GTX9_RXLOSSOFSYNC_OUT,
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    input           GTX9_GTXRXRESET_IN,
    input           GTX9_MGTREFCLKRX_IN,
    input           GTX9_PLLRXRESET_IN,
    output          GTX9_RXPLLLKDET_OUT,
    output          GTX9_RXRESETDONE_OUT,
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    output          GTX9_RXVALID_OUT,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           GTX9_RXPOLARITY_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [64:0]  GTX9_SEED_IN,
    input   [64:0]  GTX9_RXSEED,
    output          GTX9_TXOUTCLK_OUT,
    input           GTX9_TXRESET_IN,
    input           GTX9_TXUSRCLK2_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GTX9_TXN_OUT,
    output          GTX9_TXP_OUT,
    input           gtx9_force_error,
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    input           GTX9_TXDLYALIGNDISABLE_IN,
    input           GTX9_TXDLYALIGNMONENB_IN,
    output  [7:0]   GTX9_TXDLYALIGNMONITOR_OUT,
    input           GTX9_TXDLYALIGNRESET_IN,
    input           GTX9_TXENPMAPHASEALIGN_IN,
    input           GTX9_TXPMASETPHASE_IN,
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    input           GTX9_GTXTXRESET_IN,
    output          GTX9_TXRESETDONE_OUT,

    //_________________________________________________________________________
    //_________________________________________________________________________
    //GTX10  (X0Y10)
    //---------------------- Loopback and Powerdown Ports ----------------------
//jg    input   [1:0]   GTX10_RXPOWERDOWN_IN,
//jg    input   [1:0]   GTX10_TXPOWERDOWN_IN,
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg    output  [1:0]   GTX10_RXCHARISCOMMA_OUT,
//jg    output  [1:0]   GTX10_RXDISPERR_OUT,
//jg    output  [1:0]   GTX10_RXNOTINTABLE_OUT,
    //----------------- Receive Ports - Clock Correction Ports -----------------
    output  [2:0]   GTX10_RXCLKCORCNT_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          GTX10_RXBYTEREALIGN_OUT,
    output          GTX10_RXCOMMADET_OUT,
    input           GTX10_RXENMCOMMAALIGN_IN,
    input           GTX10_RXENPCOMMAALIGN_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
//jg    output  [15:0]  GTX10_RXDATA_OUT,
    input           GTX10_RXRESET_IN,
    input           GTX10_RXUSRCLK2_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input           GTX10_RXCDRRESET_IN,
    input           GTX10_RXN_IN,
    input           GTX10_RXP_IN,
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg    output  [2:0]   GTX10_RXBUFSTATUS_OUT,
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    output  [1:0]   GTX10_RXLOSSOFSYNC_OUT,
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    input           GTX10_GTXRXRESET_IN,
    input           GTX10_MGTREFCLKRX_IN,
    input           GTX10_PLLRXRESET_IN,
    output          GTX10_RXPLLLKDET_OUT,
    output          GTX10_RXRESETDONE_OUT,
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    output          GTX10_RXVALID_OUT,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           GTX10_RXPOLARITY_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [64:0]  GTX10_SEED_IN,
    input   [64:0]  GTX10_RXSEED,
    output          GTX10_TXOUTCLK_OUT,
    input           GTX10_TXRESET_IN,
    input           GTX10_TXUSRCLK2_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GTX10_TXN_OUT,
    output          GTX10_TXP_OUT,
    input           gtx10_force_error,
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    input           GTX10_TXDLYALIGNDISABLE_IN,
    input           GTX10_TXDLYALIGNMONENB_IN,
    output  [7:0]   GTX10_TXDLYALIGNMONITOR_OUT,
    input           GTX10_TXDLYALIGNRESET_IN,
    input           GTX10_TXENPMAPHASEALIGN_IN,
    input           GTX10_TXPMASETPHASE_IN,
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    input           GTX10_GTXTXRESET_IN,
    output          GTX10_TXRESETDONE_OUT,

    //_________________________________________________________________________
    //_________________________________________________________________________
    //GTX11  (X0Y11)
    //---------------------- Loopback and Powerdown Ports ----------------------
//jg    input   [1:0]   GTX11_RXPOWERDOWN_IN,
//jg    input   [1:0]   GTX11_TXPOWERDOWN_IN,
    //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg    output  [1:0]   GTX11_RXCHARISCOMMA_OUT,
//jg    output  [1:0]   GTX11_RXDISPERR_OUT,
//jg    output  [1:0]   GTX11_RXNOTINTABLE_OUT,
    //----------------- Receive Ports - Clock Correction Ports -----------------
    output  [2:0]   GTX11_RXCLKCORCNT_OUT,
    //------------- Receive Ports - Comma Detection and Alignment --------------
    output          GTX11_RXBYTEREALIGN_OUT,
    output          GTX11_RXCOMMADET_OUT,
    input           GTX11_RXENMCOMMAALIGN_IN,
    input           GTX11_RXENPCOMMAALIGN_IN,
    //----------------- Receive Ports - RX Data Path interface -----------------
//jg    output  [15:0]  GTX11_RXDATA_OUT,
    input           GTX11_RXRESET_IN,
    input           GTX11_RXUSRCLK2_IN,
    //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    input           GTX11_RXCDRRESET_IN,
    input           GTX11_RXN_IN,
    input           GTX11_RXP_IN,
    //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg    output  [2:0]   GTX11_RXBUFSTATUS_OUT,
    //------------- Receive Ports - RX Loss-of-sync State Machine --------------
    output  [1:0]   GTX11_RXLOSSOFSYNC_OUT,
    //---------------------- Receive Ports - RX PLL Ports ----------------------
    input           GTX11_GTXRXRESET_IN,
    input           GTX11_MGTREFCLKRX_IN,
    input           GTX11_PLLRXRESET_IN,
    output          GTX11_RXPLLLKDET_OUT,
    output          GTX11_RXRESETDONE_OUT,
    //------------ Receive Ports - RX Pipe Control for PCI Express -------------
    output          GTX11_RXVALID_OUT,
    //--------------- Receive Ports - RX Polarity Control Ports ----------------
    input           GTX11_RXPOLARITY_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [64:0]  GTX11_SEED_IN,
    input   [64:0]  GTX11_RXSEED,
    output          GTX11_TXOUTCLK_OUT,
    input           GTX11_TXRESET_IN,
    input           GTX11_TXUSRCLK2_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GTX11_TXN_OUT,
    output          GTX11_TXP_OUT,
    input           gtx11_force_error,
    //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
    input           GTX11_TXDLYALIGNDISABLE_IN,
    input           GTX11_TXDLYALIGNMONENB_IN,
    output  [7:0]   GTX11_TXDLYALIGNMONITOR_OUT,
    input           GTX11_TXDLYALIGNRESET_IN,
    input           GTX11_TXENPMAPHASEALIGN_IN,
    input           GTX11_TXPMASETPHASE_IN,
    //--------------------- Transmit Ports - TX PLL Ports ----------------------
    input           GTX11_GTXTXRESET_IN,
    output          GTX11_TXRESETDONE_OUT
);

//***************************** Wire Declarations *****************************
    // ground and vcc signals
    wire           tied_to_ground_i;
    wire   [63:0]  tied_to_ground_vec_i;
    wire           tied_to_vcc_i;
    wire   [63:0]  tied_to_vcc_vec_i;
    wire   [1:0]   low2, high2;
   
//********************************* Main Body of Code**************************
    assign tied_to_ground_i             = 1'b0;
    assign tied_to_ground_vec_i         = 64'h0000000000000000;
    assign tied_to_vcc_i                = 1'b1;
    assign tied_to_vcc_vec_i            = 64'hffffffffffffffff;
    assign low2  = 2'b00;
    assign high2 = 2'b11;

//------------------------- GTX Instances  -------------------------------

//_________________________________________________________________________
//_________________________________________________________________________
//GTX0  (X0Y0)  TX9-fiber6 + RX0-fiber1[boardRX0]
    SNAP12_T20R20_GTX #
    (
        // Simulation attributes
        .GTX_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        // Share RX PLL parameter
        .GTX_TX_CLK_SOURCE           ("RXPLL"),
        // Save power parameter
        //old .GTX_POWER_SAVE              (10'b0000100100)
// new default      
        .GTX_POWER_SAVE              (10'b0000110000)
    )
    gtx0_snap12_t20r20_i
    (
        //---------------------- Loopback and Powerdown Ports ----------------------
        .RXPOWERDOWN_IN                 (low2),
        .TXPOWERDOWN_IN                 (low2),
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg        .RXCHARISCOMMA_OUT              (GTX0_RXCHARISCOMMA_OUT),
//jg        .RXCHARISK_OUT                  (GTX1_RXCHARISK_OUT),
//jg        .RXDISPERR_OUT                  (GTX0_RXDISPERR_OUT),
//jg        .RXNOTINTABLE_OUT               (GTX0_RXNOTINTABLE_OUT),
        .gtx_wait  (gtx_wait),
        .rxdv      (rxdv_snapr[0]),
        .rxcomma   (rxcomma_snapr[0]),
        .check_ok  (check_ok_snapr[0]),
        .check_bad (check_bad_snapr[0]),
        .good_byte (good_byte[0]),
        .bad_byte  (bad_byte[0]),
        .lost_byte (lost_byte[0]),
        .err_count (errcount0),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .RXCLKCORCNT_OUT                (GTX0_RXCLKCORCNT_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEREALIGN_OUT              (GTX0_RXBYTEREALIGN_OUT),
        .RXCOMMADET_OUT                 (GTX0_RXCOMMADET_OUT),
        .RXENMCOMMAALIGN_IN             (GTX0_RXENMCOMMAALIGN_IN),
        .RXENPCOMMAALIGN_IN             (GTX0_RXENPCOMMAALIGN_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA_OUT                     (),
        .RXCHARISK_OUT                  (),
        .RXRESET_IN                     (GTX0_RXRESET_IN),
        .RXUSRCLK2_IN                   (GTX0_RXUSRCLK2_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXCDRRESET_IN                  (GTX0_RXCDRRESET_IN),
        .RXN_IN                         (GTX0_RXN_IN),
        .RXP_IN                         (GTX0_RXP_IN),
        //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg        .RXBUFSTATUS_OUT                (GTX0_RXBUFSTATUS_OUT),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .RXLOSSOFSYNC_OUT               (GTX0_RXLOSSOFSYNC_OUT),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTXRXRESET_IN                  (GTX0_GTXRXRESET_IN),
        .MGTREFCLKRX_IN                 ({tied_to_ground_i , GTX0_MGTREFCLKRX_IN}),
        .PLLRXRESET_IN                  (GTX0_PLLRXRESET_IN),
        .RXPLLLKDET_OUT                 (GTX0_RXPLLLKDET_OUT),
        .RXRESETDONE_OUT                (GTX0_RXRESETDONE_OUT),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .RXVALID_OUT                    (GTX0_RXVALID_OUT),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY_IN                  (GTX0_RXPOLARITY_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .iseed                       (GTX0_SEED_IN),
        .rxseed                      (GTX0_RXSEED),
        .force_error                 (gtx0_force_error),
        .TXOUTCLK_OUT                   (GTX0_TXOUTCLK_OUT),
        .TXRESET_IN                     (GTX0_TXRESET_IN),
        .TXUSRCLK2_IN                   (GTX0_TXUSRCLK2_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .TXN_OUT                        (GTX0_TXN_OUT),
        .TXP_OUT                        (GTX0_TXP_OUT),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .TXDLYALIGNDISABLE_IN           (GTX0_TXDLYALIGNDISABLE_IN),
        .TXDLYALIGNMONENB_IN            (GTX0_TXDLYALIGNMONENB_IN),
        .TXDLYALIGNMONITOR_OUT          (GTX0_TXDLYALIGNMONITOR_OUT),
        .TXDLYALIGNRESET_IN             (GTX0_TXDLYALIGNRESET_IN),
        .TXENPMAPHASEALIGN_IN           (GTX0_TXENPMAPHASEALIGN_IN),
        .TXPMASETPHASE_IN               (GTX0_TXPMASETPHASE_IN),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTXTXRESET_IN                  (GTX0_GTXTXRESET_IN),
        .MGTREFCLKTX_IN                 ({tied_to_ground_i , GTX0_MGTREFCLKRX_IN}),
        .PLLTXRESET_IN                  (tied_to_ground_i),
        .TXPLLLKDET_OUT                 (),
        .TXRESETDONE_OUT                (GTX0_TXRESETDONE_OUT)
    );

//_________________________________________________________________________
//_________________________________________________________________________
//GTX1  (X0Y1)  TX8-fiber5 + RX1-fiber2[boardRX1]
    SNAP12_T20R20_GTX #
    (
        // Simulation attributes
        .GTX_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        // Share RX PLL parameter
        .GTX_TX_CLK_SOURCE           ("RXPLL"),
        // Save power parameter
        //old .GTX_POWER_SAVE              (10'b0000100100)
// new default        
        .GTX_POWER_SAVE              (10'b0000110000)
    )
    gtx1_snap12_t20r20_i
    (
        //---------------------- Loopback and Powerdown Ports ----------------------
        .RXPOWERDOWN_IN                 (low2),
        .TXPOWERDOWN_IN                 (low2),
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg        .RXCHARISCOMMA_OUT              (GTX1_RXCHARISCOMMA_OUT),
//jg        .RXCHARISK_OUT                  (GTX1_RXCHARISK_OUT),
//jg        .RXDISPERR_OUT                  (GTX1_RXDISPERR_OUT),
//jg        .RXNOTINTABLE_OUT               (GTX1_RXNOTINTABLE_OUT),
        .gtx_wait  (gtx_wait),
        .rxdv      (rxdv_snapr[1]),
        .rxcomma   (rxcomma_snapr[1]),
        .check_ok  (check_ok_snapr[1]),
        .check_bad (check_bad_snapr[1]),
        .good_byte (good_byte[1]),
        .bad_byte  (bad_byte[1]),
        .lost_byte (lost_byte[1]),
        .err_count (errcount1),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .RXCLKCORCNT_OUT                (GTX1_RXCLKCORCNT_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEREALIGN_OUT              (GTX1_RXBYTEREALIGN_OUT),
        .RXCOMMADET_OUT                 (GTX1_RXCOMMADET_OUT),
        .RXENMCOMMAALIGN_IN             (GTX1_RXENMCOMMAALIGN_IN),
        .RXENPCOMMAALIGN_IN             (GTX1_RXENPCOMMAALIGN_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA_OUT                     (GTXi_RXDATA_OUT),  // select just ONE gtx data to monitor...
        .RXCHARISK_OUT                  (GTXi_RXK_OUT),     // select the K that goes with it
//JGtemp        .RXDATA_OUT                     (),
//JGtemp        .RXCHARISK_OUT                  (),
        .RXRESET_IN                     (GTX1_RXRESET_IN),
        .RXUSRCLK2_IN                   (GTX1_RXUSRCLK2_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXCDRRESET_IN                  (GTX1_RXCDRRESET_IN),
        .RXN_IN                         (GTX1_RXN_IN),
        .RXP_IN                         (GTX1_RXP_IN),
        //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg        .RXBUFSTATUS_OUT                (GTX1_RXBUFSTATUS_OUT),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .RXLOSSOFSYNC_OUT               (GTX1_RXLOSSOFSYNC_OUT),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTXRXRESET_IN                  (GTX1_GTXRXRESET_IN),
        .MGTREFCLKRX_IN                 ({tied_to_ground_i , GTX1_MGTREFCLKRX_IN}),
        .PLLRXRESET_IN                  (GTX1_PLLRXRESET_IN),
        .RXPLLLKDET_OUT                 (GTX1_RXPLLLKDET_OUT),
        .RXRESETDONE_OUT                (GTX1_RXRESETDONE_OUT),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .RXVALID_OUT                    (GTX1_RXVALID_OUT),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY_IN                  (GTX1_RXPOLARITY_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .iseed                       (GTX1_SEED_IN),
        .rxseed                      (GTX1_RXSEED),
        .force_error                 (gtx1_force_error),
        .TXOUTCLK_OUT                   (GTX1_TXOUTCLK_OUT),
        .TXRESET_IN                     (GTX1_TXRESET_IN),
        .TXUSRCLK2_IN                   (GTX1_TXUSRCLK2_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .TXN_OUT                        (GTX1_TXN_OUT),
        .TXP_OUT                        (GTX1_TXP_OUT),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .TXDLYALIGNDISABLE_IN           (GTX1_TXDLYALIGNDISABLE_IN),
        .TXDLYALIGNMONENB_IN            (GTX1_TXDLYALIGNMONENB_IN),
        .TXDLYALIGNMONITOR_OUT          (GTX1_TXDLYALIGNMONITOR_OUT),
        .TXDLYALIGNRESET_IN             (GTX1_TXDLYALIGNRESET_IN),
        .TXENPMAPHASEALIGN_IN           (GTX1_TXENPMAPHASEALIGN_IN),
        .TXPMASETPHASE_IN               (GTX1_TXPMASETPHASE_IN),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTXTXRESET_IN                  (GTX1_GTXTXRESET_IN),
        .MGTREFCLKTX_IN                 ({tied_to_ground_i , GTX1_MGTREFCLKRX_IN}),
        .PLLTXRESET_IN                  (tied_to_ground_i),
        .TXPLLLKDET_OUT                 (),
        .TXRESETDONE_OUT                (GTX1_TXRESETDONE_OUT)
    );

//_________________________________________________________________________
//_________________________________________________________________________
//GTX2  (X0Y2)  TX7-fiber12 + RX2-fiber3[boardRX2]
    SNAP12_T20R20_GTX #
    (
        // Simulation attributes
        .GTX_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        // Share RX PLL parameter
        .GTX_TX_CLK_SOURCE           ("RXPLL"),
        // Save power parameter
        // old .GTX_POWER_SAVE              (10'b0000100100)
// new default        
        .GTX_POWER_SAVE              (10'b0000110000)
    )
    gtx2_snap12_t20r20_i
    (
        //---------------------- Loopback and Powerdown Ports ----------------------
        .RXPOWERDOWN_IN                 (low2),
        .TXPOWERDOWN_IN                 (low2),
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg        .RXCHARISCOMMA_OUT              (GTX2_RXCHARISCOMMA_OUT),
//jg        .RXCHARISK_OUT                  (GTX2_RXCHARISK_OUT),
//jg        .RXDISPERR_OUT                  (GTX2_RXDISPERR_OUT),
//jg        .RXNOTINTABLE_OUT               (GTX2_RXNOTINTABLE_OUT),
        .gtx_wait  (gtx_wait),
        .rxdv      (rxdv_snapr[2]),
        .rxcomma   (rxcomma_snapr[2]),
        .check_ok  (check_ok_snapr[2]),
        .check_bad (check_bad_snapr[2]),
        .good_byte (good_byte[2]),
        .bad_byte  (bad_byte[2]),
        .lost_byte (lost_byte[2]),
        .err_count (errcount2),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .RXCLKCORCNT_OUT                (GTX2_RXCLKCORCNT_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEREALIGN_OUT              (GTX2_RXBYTEREALIGN_OUT),
        .RXCOMMADET_OUT                 (GTX2_RXCOMMADET_OUT),
        .RXENMCOMMAALIGN_IN             (GTX2_RXENMCOMMAALIGN_IN),
        .RXENPCOMMAALIGN_IN             (GTX2_RXENPCOMMAALIGN_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA_OUT                     (),
        .RXCHARISK_OUT                  (),
        .RXRESET_IN                     (GTX2_RXRESET_IN),
        .RXUSRCLK2_IN                   (GTX2_RXUSRCLK2_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXCDRRESET_IN                  (GTX2_RXCDRRESET_IN),
        .RXN_IN                         (GTX2_RXN_IN),
        .RXP_IN                         (GTX2_RXP_IN),
        //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg        .RXBUFSTATUS_OUT                (GTX2_RXBUFSTATUS_OUT),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .RXLOSSOFSYNC_OUT               (GTX2_RXLOSSOFSYNC_OUT),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTXRXRESET_IN                  (GTX2_GTXRXRESET_IN),
        .MGTREFCLKRX_IN                 ({tied_to_ground_i , GTX2_MGTREFCLKRX_IN}),
        .PLLRXRESET_IN                  (GTX2_PLLRXRESET_IN),
        .RXPLLLKDET_OUT                 (GTX2_RXPLLLKDET_OUT),
        .RXRESETDONE_OUT                (GTX2_RXRESETDONE_OUT),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .RXVALID_OUT                    (GTX2_RXVALID_OUT),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY_IN                  (GTX2_RXPOLARITY_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .iseed                       (GTX2_SEED_IN),
        .rxseed                      (GTX2_RXSEED),
        .force_error                 (gtx2_force_error),
        .TXOUTCLK_OUT                   (GTX2_TXOUTCLK_OUT),
        .TXRESET_IN                     (GTX2_TXRESET_IN),
        .TXUSRCLK2_IN                   (GTX2_TXUSRCLK2_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .TXN_OUT                        (GTX2_TXN_OUT),
        .TXP_OUT                        (GTX2_TXP_OUT),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .TXDLYALIGNDISABLE_IN           (GTX2_TXDLYALIGNDISABLE_IN),
        .TXDLYALIGNMONENB_IN            (GTX2_TXDLYALIGNMONENB_IN),
        .TXDLYALIGNMONITOR_OUT          (GTX2_TXDLYALIGNMONITOR_OUT),
        .TXDLYALIGNRESET_IN             (GTX2_TXDLYALIGNRESET_IN),
        .TXENPMAPHASEALIGN_IN           (GTX2_TXENPMAPHASEALIGN_IN),
        .TXPMASETPHASE_IN               (GTX2_TXPMASETPHASE_IN),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTXTXRESET_IN                  (GTX2_GTXTXRESET_IN),
        .MGTREFCLKTX_IN                 ({tied_to_ground_i , GTX2_MGTREFCLKRX_IN}),
        .PLLTXRESET_IN                  (tied_to_ground_i),
        .TXPLLLKDET_OUT                 (),
        .TXRESETDONE_OUT                (GTX2_TXRESETDONE_OUT)
    );

//_________________________________________________________________________
//_________________________________________________________________________
//GTX3  (X0Y3)  TX0-fiber1 + RX3-fiber4[boardRX3]
    SNAP12_T20R20_GTX #
    (
        // Simulation attributes
        .GTX_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        // Share RX PLL parameter
        .GTX_TX_CLK_SOURCE           ("RXPLL"),
        // Save power parameter
        //old  .GTX_POWER_SAVE              (10'b0000100100)
// new default        
        .GTX_POWER_SAVE              (10'b0000110000)
    )
    gtx3_snap12_t20r20_i
    (
        //---------------------- Loopback and Powerdown Ports ----------------------
        .RXPOWERDOWN_IN                 (low2),
        .TXPOWERDOWN_IN                 (low2),
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg        .RXCHARISCOMMA_OUT              (GTX3_RXCHARISCOMMA_OUT),
//jg        .RXCHARISK_OUT                  (GTX3_RXCHARISK_OUT),
//jg        .RXDISPERR_OUT                  (GTX3_RXDISPERR_OUT),
//jg        .RXNOTINTABLE_OUT               (GTX3_RXNOTINTABLE_OUT),
        .gtx_wait  (gtx_wait),
        .rxdv      (rxdv_snapr[3]),
        .rxcomma   (rxcomma_snapr[3]),
        .check_ok  (check_ok_snapr[3]),
        .check_bad (check_bad_snapr[3]),
        .good_byte (good_byte[3]),
        .bad_byte  (bad_byte[3]),
        .lost_byte (lost_byte[3]),
        .err_count (errcount3),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .RXCLKCORCNT_OUT                (GTX3_RXCLKCORCNT_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEREALIGN_OUT              (GTX3_RXBYTEREALIGN_OUT),
        .RXCOMMADET_OUT                 (GTX3_RXCOMMADET_OUT),
        .RXENMCOMMAALIGN_IN             (GTX3_RXENMCOMMAALIGN_IN),
        .RXENPCOMMAALIGN_IN             (GTX3_RXENPCOMMAALIGN_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA_OUT                     (),
        .RXCHARISK_OUT                  (),
        .RXRESET_IN                     (GTX3_RXRESET_IN),
        .RXUSRCLK2_IN                   (GTX3_RXUSRCLK2_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXCDRRESET_IN                  (GTX3_RXCDRRESET_IN),
        .RXN_IN                         (GTX3_RXN_IN),
        .RXP_IN                         (GTX3_RXP_IN),
        //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg        .RXBUFSTATUS_OUT                (GTX3_RXBUFSTATUS_OUT),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .RXLOSSOFSYNC_OUT               (GTX3_RXLOSSOFSYNC_OUT),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTXRXRESET_IN                  (GTX3_GTXRXRESET_IN),
        .MGTREFCLKRX_IN                 ({tied_to_ground_i , GTX3_MGTREFCLKRX_IN}),
        .PLLRXRESET_IN                  (GTX3_PLLRXRESET_IN),
        .RXPLLLKDET_OUT                 (GTX3_RXPLLLKDET_OUT),
        .RXRESETDONE_OUT                (GTX3_RXRESETDONE_OUT),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .RXVALID_OUT                    (GTX3_RXVALID_OUT),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY_IN                  (GTX3_RXPOLARITY_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .iseed                       (GTX3_SEED_IN),
        .rxseed                      (GTX3_RXSEED),
        .force_error                 (gtx3_force_error),
        .TXOUTCLK_OUT                   (GTX3_TXOUTCLK_OUT),
        .TXRESET_IN                     (GTX3_TXRESET_IN),
        .TXUSRCLK2_IN                   (GTX3_TXUSRCLK2_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .TXN_OUT                        (GTX3_TXN_OUT),
        .TXP_OUT                        (GTX3_TXP_OUT),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .TXDLYALIGNDISABLE_IN           (GTX3_TXDLYALIGNDISABLE_IN),
        .TXDLYALIGNMONENB_IN            (GTX3_TXDLYALIGNMONENB_IN),
        .TXDLYALIGNMONITOR_OUT          (GTX3_TXDLYALIGNMONITOR_OUT),
        .TXDLYALIGNRESET_IN             (GTX3_TXDLYALIGNRESET_IN),
        .TXENPMAPHASEALIGN_IN           (GTX3_TXENPMAPHASEALIGN_IN),
        .TXPMASETPHASE_IN               (GTX3_TXPMASETPHASE_IN),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTXTXRESET_IN                  (GTX3_GTXTXRESET_IN),
        .MGTREFCLKTX_IN                 ({tied_to_ground_i , GTX3_MGTREFCLKRX_IN}),
        .PLLTXRESET_IN                  (tied_to_ground_i),
        .TXPLLLKDET_OUT                 (),
        .TXRESETDONE_OUT                (GTX3_TXRESETDONE_OUT)
    );

//_________________________________________________________________________
//_________________________________________________________________________
//GTX4  (X0Y4)  TX1-fiber2 + GemRX0-fiber5[boardRX4]
    SNAP12_T20R20_GTX #
    (
        // Simulation attributes
        .GTX_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        // Share RX PLL parameter
        .GTX_TX_CLK_SOURCE           ("RXPLL"),
        // Save power parameter
        //old  .GTX_POWER_SAVE              (10'b0000100100)
// new default    
        .GTX_POWER_SAVE              (10'b0000110000)
    )
    gtx4_snap12_t20r20_i
    (
        //---------------------- Loopback and Powerdown Ports ----------------------
        .RXPOWERDOWN_IN                 (low2),
        .TXPOWERDOWN_IN                 (low2),
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg        .RXCHARISCOMMA_OUT              (GTX4_RXCHARISCOMMA_OUT),
//jg        .RXCHARISK_OUT                  (GTX4_RXCHARISK_OUT),
//jg        .RXDISPERR_OUT                  (GTX4_RXDISPERR_OUT),
//jg        .RXNOTINTABLE_OUT               (GTX4_RXNOTINTABLE_OUT),
        .gtx_wait  (gtx_wait),  // this TX goes to a different active RX, be careful!
        .rxdv      (rxdv_snapr[8]),   //JG, From here down is New!
        .rxcomma   (rxcomma_snapr[8]),
        .check_ok  (check_ok_snapr[8]),
        .check_bad (check_bad_snapr[8]),
        .good_byte (good_byte[8]),
        .bad_byte  (bad_byte[8]),
        .lost_byte (lost_byte[8]),
        .err_count (errcount8),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .RXCLKCORCNT_OUT                (GTX4_RXCLKCORCNT_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEREALIGN_OUT              (GTX4_RXBYTEREALIGN_OUT),
        .RXCOMMADET_OUT                 (GTX4_RXCOMMADET_OUT),
        .RXENMCOMMAALIGN_IN             (GTX4_RXENMCOMMAALIGN_IN),
        .RXENPCOMMAALIGN_IN             (GTX4_RXENPCOMMAALIGN_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA_OUT                     (),
        .RXCHARISK_OUT                  (),
        .RXRESET_IN                     (GTX4_RXRESET_IN),
        .RXUSRCLK2_IN                   (GTX4_RXUSRCLK2_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXCDRRESET_IN                  (GTX4_RXCDRRESET_IN),
        .RXN_IN                         (GTX4_RXN_IN),
        .RXP_IN                         (GTX4_RXP_IN),
        //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg        .RXBUFSTATUS_OUT                (GTX4_RXBUFSTATUS_OUT),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .RXLOSSOFSYNC_OUT               (GTX4_RXLOSSOFSYNC_OUT),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTXRXRESET_IN                  (GTX4_GTXRXRESET_IN),
        .MGTREFCLKRX_IN                 ({tied_to_ground_i , GTX4_MGTREFCLKRX_IN}),
        .PLLRXRESET_IN                  (GTX4_PLLRXRESET_IN),
        .RXPLLLKDET_OUT                 (GTX4_RXPLLLKDET_OUT),
        .RXRESETDONE_OUT                (GTX4_RXRESETDONE_OUT),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .RXVALID_OUT                    (GTX4_RXVALID_OUT),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY_IN                  (GTX4_RXPOLARITY_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .iseed                       (GTX4_SEED_IN),
        .rxseed                      (GTX4_RXSEED),
        .force_error                 (gtx4_force_error),
        .TXOUTCLK_OUT                   (GTX4_TXOUTCLK_OUT),
        .TXRESET_IN                     (GTX4_TXRESET_IN),
        .TXUSRCLK2_IN                   (GTX4_TXUSRCLK2_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .TXN_OUT                        (GTX4_TXN_OUT),
        .TXP_OUT                        (GTX4_TXP_OUT),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .TXDLYALIGNDISABLE_IN           (GTX4_TXDLYALIGNDISABLE_IN),
        .TXDLYALIGNMONENB_IN            (GTX4_TXDLYALIGNMONENB_IN),
        .TXDLYALIGNMONITOR_OUT          (GTX4_TXDLYALIGNMONITOR_OUT),
        .TXDLYALIGNRESET_IN             (GTX4_TXDLYALIGNRESET_IN),
        .TXENPMAPHASEALIGN_IN           (GTX4_TXENPMAPHASEALIGN_IN),
        .TXPMASETPHASE_IN               (GTX4_TXPMASETPHASE_IN),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTXTXRESET_IN                  (GTX4_GTXTXRESET_IN),
        .MGTREFCLKTX_IN                 ({tied_to_ground_i , GTX4_MGTREFCLKRX_IN}),
        .PLLTXRESET_IN                  (tied_to_ground_i),
        .TXPLLLKDET_OUT                 (),
        .TXRESETDONE_OUT                (GTX4_TXRESETDONE_OUT)
    );

//_________________________________________________________________________
//_________________________________________________________________________
//GTX5  (X0Y5)  TX11-fiber8 or GemRX1-fiber6[boardRX5]
    SNAP12_T20R20_GTX #
    (
        // Simulation attributes
        .GTX_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        // Share RX PLL parameter
        .GTX_TX_CLK_SOURCE           ("RXPLL"),
        // Save power parameter
        //old .GTX_POWER_SAVE              (10'b0000100100)
// new default       
        .GTX_POWER_SAVE              (10'b0000110000)
    )
    gtx5_snap12_t20r20_i
    (
        //---------------------- Loopback and Powerdown Ports ----------------------
        .RXPOWERDOWN_IN                 (low2),
        .TXPOWERDOWN_IN                 (low2),
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg        .RXCHARISCOMMA_OUT              (GTX5_RXCHARISCOMMA_OUT),
//jg        .RXCHARISK_OUT                  (GTX5_RXCHARISK_OUT),
//jg        .RXDISPERR_OUT                  (GTX5_RXDISPERR_OUT),
//jg        .RXNOTINTABLE_OUT               (GTX5_RXNOTINTABLE_OUT),
        .gtx_wait  (gtx_wait),   //JG, All New!
        .rxdv      (rxdv_snapr[9]),
        .rxcomma   (rxcomma_snapr[9]),
        .check_ok  (check_ok_snapr[9]),
        .check_bad (check_bad_snapr[9]),
        .good_byte (good_byte[9]),
        .bad_byte  (bad_byte[9]),
        .lost_byte (lost_byte[9]),
        .err_count (errcount9),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .RXCLKCORCNT_OUT                (GTX5_RXCLKCORCNT_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEREALIGN_OUT              (GTX5_RXBYTEREALIGN_OUT),
        .RXCOMMADET_OUT                 (GTX5_RXCOMMADET_OUT),
        .RXENMCOMMAALIGN_IN             (GTX5_RXENMCOMMAALIGN_IN),
        .RXENPCOMMAALIGN_IN             (GTX5_RXENPCOMMAALIGN_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA_OUT                     (),
        .RXCHARISK_OUT                  (),
        .RXRESET_IN                     (GTX5_RXRESET_IN),
        .RXUSRCLK2_IN                   (GTX5_RXUSRCLK2_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXCDRRESET_IN                  (GTX5_RXCDRRESET_IN),
        .RXN_IN                         (GTX5_RXN_IN),
        .RXP_IN                         (GTX5_RXP_IN),
        //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg        .RXBUFSTATUS_OUT                (GTX5_RXBUFSTATUS_OUT),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .RXLOSSOFSYNC_OUT               (GTX5_RXLOSSOFSYNC_OUT),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTXRXRESET_IN                  (GTX5_GTXRXRESET_IN),
        .MGTREFCLKRX_IN                 ({tied_to_ground_i , GTX5_MGTREFCLKRX_IN}),
        .PLLRXRESET_IN                  (GTX5_PLLRXRESET_IN),
        .RXPLLLKDET_OUT                 (GTX5_RXPLLLKDET_OUT),
        .RXRESETDONE_OUT                (GTX5_RXRESETDONE_OUT),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .RXVALID_OUT                    (GTX5_RXVALID_OUT),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY_IN                  (GTX5_RXPOLARITY_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .iseed                       (GTX5_SEED_IN),
        .rxseed                      (GTX5_RXSEED),
        .force_error                 (gtx5_force_error),
        .TXOUTCLK_OUT                   (GTX5_TXOUTCLK_OUT),
        .TXRESET_IN                     (GTX5_TXRESET_IN),
        .TXUSRCLK2_IN                   (GTX5_TXUSRCLK2_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .TXN_OUT                        (GTX5_TXN_OUT),
        .TXP_OUT                        (GTX5_TXP_OUT),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .TXDLYALIGNDISABLE_IN           (GTX5_TXDLYALIGNDISABLE_IN),
        .TXDLYALIGNMONENB_IN            (GTX5_TXDLYALIGNMONENB_IN),
        .TXDLYALIGNMONITOR_OUT          (GTX5_TXDLYALIGNMONITOR_OUT),
        .TXDLYALIGNRESET_IN             (GTX5_TXDLYALIGNRESET_IN),
        .TXENPMAPHASEALIGN_IN           (GTX5_TXENPMAPHASEALIGN_IN),
        .TXPMASETPHASE_IN               (GTX5_TXPMASETPHASE_IN),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTXTXRESET_IN                  (GTX5_GTXTXRESET_IN),
        .MGTREFCLKTX_IN                 ({tied_to_ground_i , GTX5_MGTREFCLKRX_IN}),
        .PLLTXRESET_IN                  (tied_to_ground_i),
        .TXPLLLKDET_OUT                 (),
        .TXRESETDONE_OUT                (GTX5_TXRESETDONE_OUT)
    );

//_________________________________________________________________________
//_________________________________________________________________________
//GTX6  (X0Y6)  TX10-fiber7 + GemRX2-fiber7[boardRX6]
    SNAP12_T20R20_GTX #
    (
        // Simulation attributes
        .GTX_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        // Share RX PLL parameter
        .GTX_TX_CLK_SOURCE           ("RXPLL"),
        // Save power parameter
        //old  .GTX_POWER_SAVE              (10'b0000100100)
// new default      
        .GTX_POWER_SAVE              (10'b0000110000)
    )
    gtx6_snap12_t20r20_i
    (
        //---------------------- Loopback and Powerdown Ports ----------------------
        .RXPOWERDOWN_IN                 (low2),
        .TXPOWERDOWN_IN                 (low2),
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg        .RXCHARISCOMMA_OUT              (GTX6_RXCHARISCOMMA_OUT),
//jg        .RXCHARISK_OUT                  (GTX6_RXCHARISK_OUT),
//jg        .RXDISPERR_OUT                  (GTX6_RXDISPERR_OUT),
//jg        .RXNOTINTABLE_OUT               (GTX6_RXNOTINTABLE_OUT),
        .gtx_wait  (gtx_wait),   //JG, All New!
        .rxdv      (rxdv_snapr[10]),
        .rxcomma   (rxcomma_snapr[10]),
        .check_ok  (check_ok_snapr[10]),
        .check_bad (check_bad_snapr[10]),
        .good_byte (good_byte[10]),
        .bad_byte  (bad_byte[10]),
        .lost_byte (lost_byte[10]),
        .err_count (errcount10),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .RXCLKCORCNT_OUT                (GTX6_RXCLKCORCNT_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEREALIGN_OUT              (GTX6_RXBYTEREALIGN_OUT),
        .RXCOMMADET_OUT                 (GTX6_RXCOMMADET_OUT),
        .RXENMCOMMAALIGN_IN             (GTX6_RXENMCOMMAALIGN_IN),
        .RXENPCOMMAALIGN_IN             (GTX6_RXENPCOMMAALIGN_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA_OUT                     (),
        .RXCHARISK_OUT                  (),
        .RXRESET_IN                     (GTX6_RXRESET_IN),
        .RXUSRCLK2_IN                   (GTX6_RXUSRCLK2_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXCDRRESET_IN                  (GTX6_RXCDRRESET_IN),
        .RXN_IN                         (GTX6_RXN_IN),
        .RXP_IN                         (GTX6_RXP_IN),
        //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg        .RXBUFSTATUS_OUT                (GTX6_RXBUFSTATUS_OUT),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .RXLOSSOFSYNC_OUT               (GTX6_RXLOSSOFSYNC_OUT),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTXRXRESET_IN                  (GTX6_GTXRXRESET_IN),
        .MGTREFCLKRX_IN                 ({tied_to_ground_i , GTX6_MGTREFCLKRX_IN}),
        .PLLRXRESET_IN                  (GTX6_PLLRXRESET_IN),
        .RXPLLLKDET_OUT                 (GTX6_RXPLLLKDET_OUT),
        .RXRESETDONE_OUT                (GTX6_RXRESETDONE_OUT),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .RXVALID_OUT                    (GTX6_RXVALID_OUT),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY_IN                  (GTX6_RXPOLARITY_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .iseed                       (GTX6_SEED_IN),
        .rxseed                      (GTX6_RXSEED),
        .force_error                 (gtx6_force_error),
        .TXOUTCLK_OUT                   (GTX6_TXOUTCLK_OUT),
        .TXRESET_IN                     (GTX6_TXRESET_IN),
        .TXUSRCLK2_IN                   (GTX6_TXUSRCLK2_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .TXN_OUT                        (GTX6_TXN_OUT),
        .TXP_OUT                        (GTX6_TXP_OUT),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .TXDLYALIGNDISABLE_IN           (GTX6_TXDLYALIGNDISABLE_IN),
        .TXDLYALIGNMONENB_IN            (GTX6_TXDLYALIGNMONENB_IN),
        .TXDLYALIGNMONITOR_OUT          (GTX6_TXDLYALIGNMONITOR_OUT),
        .TXDLYALIGNRESET_IN             (GTX6_TXDLYALIGNRESET_IN),
        .TXENPMAPHASEALIGN_IN           (GTX6_TXENPMAPHASEALIGN_IN),
        .TXPMASETPHASE_IN               (GTX6_TXPMASETPHASE_IN),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTXTXRESET_IN                  (GTX6_GTXTXRESET_IN),
        .MGTREFCLKTX_IN                 ({tied_to_ground_i , GTX6_MGTREFCLKRX_IN}),
        .PLLTXRESET_IN                  (tied_to_ground_i),
        .TXPLLLKDET_OUT                 (),
        .TXRESETDONE_OUT                (GTX6_TXRESETDONE_OUT)
    );

//_________________________________________________________________________
//_________________________________________________________________________
//GTX7  (X0Y7)  TX2-fiber3 + GemRX3-fiber8[boardRX7]
    SNAP12_T20R20_GTX #
    (
        // Simulation attributes
        .GTX_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        // Share RX PLL parameter
        .GTX_TX_CLK_SOURCE           ("RXPLL"),
        // Save power parameter
        // old .GTX_POWER_SAVE              (10'b0000100100)
// new default        
        .GTX_POWER_SAVE              (10'b0000110000)
    )
    gtx7_snap12_t20r20_i
    (
        //---------------------- Loopback and Powerdown Ports ----------------------
        .RXPOWERDOWN_IN                 (low2),
        .TXPOWERDOWN_IN                 (low2),
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg        .RXCHARISCOMMA_OUT              (GTX7_RXCHARISCOMMA_OUT),
//jg        .RXCHARISK_OUT                  (GTX7_RXCHARISK_OUT),
//jg        .RXDISPERR_OUT                  (GTX7_RXDISPERR_OUT),
//jg        .RXNOTINTABLE_OUT               (GTX7_RXNOTINTABLE_OUT),
        .gtx_wait  (gtx_wait),  // this TX goes to a different active RX, be careful!
        .rxdv      (rxdv_snapr[11]),   //JG, From here down is New!
        .rxcomma   (rxcomma_snapr[11]),
        .check_ok  (check_ok_snapr[11]),
        .check_bad (check_bad_snapr[11]),
        .good_byte (good_byte[11]),
        .bad_byte  (bad_byte[11]),
        .lost_byte (lost_byte[11]),
        .err_count (errcount11),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .RXCLKCORCNT_OUT                (GTX7_RXCLKCORCNT_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEREALIGN_OUT              (GTX7_RXBYTEREALIGN_OUT),
        .RXCOMMADET_OUT                 (GTX7_RXCOMMADET_OUT),
        .RXENMCOMMAALIGN_IN             (GTX7_RXENMCOMMAALIGN_IN),
        .RXENPCOMMAALIGN_IN             (GTX7_RXENPCOMMAALIGN_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA_OUT                     (),
        .RXCHARISK_OUT                  (),
        .RXRESET_IN                     (GTX7_RXRESET_IN),
        .RXUSRCLK2_IN                   (GTX7_RXUSRCLK2_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXCDRRESET_IN                  (GTX7_RXCDRRESET_IN),
        .RXN_IN                         (GTX7_RXN_IN),
        .RXP_IN                         (GTX7_RXP_IN),
        //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg        .RXBUFSTATUS_OUT                (GTX7_RXBUFSTATUS_OUT),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .RXLOSSOFSYNC_OUT               (GTX7_RXLOSSOFSYNC_OUT),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTXRXRESET_IN                  (GTX7_GTXRXRESET_IN),
        .MGTREFCLKRX_IN                 ({tied_to_ground_i , GTX7_MGTREFCLKRX_IN}),
        .PLLRXRESET_IN                  (GTX7_PLLRXRESET_IN),
        .RXPLLLKDET_OUT                 (GTX7_RXPLLLKDET_OUT),
        .RXRESETDONE_OUT                (GTX7_RXRESETDONE_OUT),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .RXVALID_OUT                    (GTX7_RXVALID_OUT),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY_IN                  (GTX7_RXPOLARITY_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .iseed                       (GTX7_SEED_IN),
        .rxseed                      (GTX7_RXSEED),
        .force_error                 (gtx7_force_error),
        .TXOUTCLK_OUT                   (GTX7_TXOUTCLK_OUT),
        .TXRESET_IN                     (GTX7_TXRESET_IN),
        .TXUSRCLK2_IN                   (GTX7_TXUSRCLK2_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .TXN_OUT                        (GTX7_TXN_OUT),
        .TXP_OUT                        (GTX7_TXP_OUT),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .TXDLYALIGNDISABLE_IN           (GTX7_TXDLYALIGNDISABLE_IN),
        .TXDLYALIGNMONENB_IN            (GTX7_TXDLYALIGNMONENB_IN),
        .TXDLYALIGNMONITOR_OUT          (GTX7_TXDLYALIGNMONITOR_OUT),
        .TXDLYALIGNRESET_IN             (GTX7_TXDLYALIGNRESET_IN),
        .TXENPMAPHASEALIGN_IN           (GTX7_TXENPMAPHASEALIGN_IN),
        .TXPMASETPHASE_IN               (GTX7_TXPMASETPHASE_IN),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTXTXRESET_IN                  (GTX7_GTXTXRESET_IN),
        .MGTREFCLKTX_IN                 ({tied_to_ground_i , GTX7_MGTREFCLKRX_IN}),
        .PLLTXRESET_IN                  (tied_to_ground_i),
        .TXPLLLKDET_OUT                 (),
        .TXRESETDONE_OUT                (GTX7_TXRESETDONE_OUT)
    );

//_________________________________________________________________________
//_________________________________________________________________________
//GTX8  (X0Y8)  TX3-fiber4 + RX4-fiber9[boardRX8]
    SNAP12_T20R20_GTX #
    (
        // Simulation attributes
        .GTX_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        // Share RX PLL parameter
        .GTX_TX_CLK_SOURCE           ("RXPLL"),
        // Save power parameter
        // .GTX_POWER_SAVE              (10'b0000100100)
// new default        
        .GTX_POWER_SAVE              (10'b0000110000)
    )
    gtx8_snap12_t20r20_i
    (
        //---------------------- Loopback and Powerdown Ports ----------------------
        .RXPOWERDOWN_IN                 (low2),
        .TXPOWERDOWN_IN                 (low2),
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg        .RXCHARISCOMMA_OUT              (GTX8_RXCHARISCOMMA_OUT),
//jg        .RXCHARISK_OUT                  (GTX8_RXCHARISK_OUT),
//jg        .RXDISPERR_OUT                  (GTX8_RXDISPERR_OUT),
//jg        .RXNOTINTABLE_OUT               (GTX8_RXNOTINTABLE_OUT),
        .gtx_wait  (gtx_wait),
        .rxdv      (rxdv_snapr[4]),
        .rxcomma   (rxcomma_snapr[4]),
        .check_ok  (check_ok_snapr[4]),
        .check_bad (check_bad_snapr[4]),
        .good_byte (good_byte[4]),
        .bad_byte  (bad_byte[4]),
        .lost_byte (lost_byte[4]),
        .err_count (errcount4),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .RXCLKCORCNT_OUT                (GTX8_RXCLKCORCNT_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEREALIGN_OUT              (GTX8_RXBYTEREALIGN_OUT),
        .RXCOMMADET_OUT                 (GTX8_RXCOMMADET_OUT),
        .RXENMCOMMAALIGN_IN             (GTX8_RXENMCOMMAALIGN_IN),
        .RXENPCOMMAALIGN_IN             (GTX8_RXENPCOMMAALIGN_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA_OUT                     (),
        .RXCHARISK_OUT                  (),
        .RXRESET_IN                     (GTX8_RXRESET_IN),
        .RXUSRCLK2_IN                   (GTX8_RXUSRCLK2_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXCDRRESET_IN                  (GTX8_RXCDRRESET_IN),
        .RXN_IN                         (GTX8_RXN_IN),
        .RXP_IN                         (GTX8_RXP_IN),
        //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg        .RXBUFSTATUS_OUT                (GTX8_RXBUFSTATUS_OUT),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .RXLOSSOFSYNC_OUT               (GTX8_RXLOSSOFSYNC_OUT),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTXRXRESET_IN                  (GTX8_GTXRXRESET_IN),
        .MGTREFCLKRX_IN                 ({tied_to_ground_i , GTX8_MGTREFCLKRX_IN}),
        .PLLRXRESET_IN                  (GTX8_PLLRXRESET_IN),
        .RXPLLLKDET_OUT                 (GTX8_RXPLLLKDET_OUT),
        .RXRESETDONE_OUT                (GTX8_RXRESETDONE_OUT),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .RXVALID_OUT                    (GTX8_RXVALID_OUT),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY_IN                  (GTX8_RXPOLARITY_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .iseed                       (GTX8_SEED_IN),
        .rxseed                      (GTX8_RXSEED),
        .force_error                 (gtx8_force_error),
        .TXOUTCLK_OUT                   (GTX8_TXOUTCLK_OUT),
        .TXRESET_IN                     (GTX8_TXRESET_IN),
        .TXUSRCLK2_IN                   (GTX8_TXUSRCLK2_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .TXN_OUT                        (GTX8_TXN_OUT),
        .TXP_OUT                        (GTX8_TXP_OUT),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .TXDLYALIGNDISABLE_IN           (GTX8_TXDLYALIGNDISABLE_IN),
        .TXDLYALIGNMONENB_IN            (GTX8_TXDLYALIGNMONENB_IN),
        .TXDLYALIGNMONITOR_OUT          (GTX8_TXDLYALIGNMONITOR_OUT),
        .TXDLYALIGNRESET_IN             (GTX8_TXDLYALIGNRESET_IN),
        .TXENPMAPHASEALIGN_IN           (GTX8_TXENPMAPHASEALIGN_IN),
        .TXPMASETPHASE_IN               (GTX8_TXPMASETPHASE_IN),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTXTXRESET_IN                  (GTX8_GTXTXRESET_IN),
        .MGTREFCLKTX_IN                 ({tied_to_ground_i , GTX8_MGTREFCLKRX_IN}),
        .PLLTXRESET_IN                  (tied_to_ground_i),
        .TXPLLLKDET_OUT                 (),
        .TXRESETDONE_OUT                (GTX8_TXRESETDONE_OUT)
    );

//_________________________________________________________________________
//_________________________________________________________________________
//GTX9  (X0Y9)  TX4-fiber9 + RX5-fiber10[boardRX9]
    SNAP12_T20R20_GTX #
    (
        // Simulation attributes
        .GTX_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        // Share RX PLL parameter
        .GTX_TX_CLK_SOURCE           ("RXPLL"),
        // Save power parameter
        //old  .GTX_POWER_SAVE              (10'b0000100100)
// new default     
        .GTX_POWER_SAVE              (10'b0000110000)
    )
    gtx9_snap12_t20r20_i
    (
        //---------------------- Loopback and Powerdown Ports ----------------------
        .RXPOWERDOWN_IN                 (low2),
        .TXPOWERDOWN_IN                 (low2),
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg        .RXCHARISCOMMA_OUT              (GTX9_RXCHARISCOMMA_OUT),
//jg        .RXCHARISK_OUT                  (GTX9_RXCHARISK_OUT),
//jg        .RXDISPERR_OUT                  (GTX9_RXDISPERR_OUT),
//jg        .RXNOTINTABLE_OUT               (GTX9_RXNOTINTABLE_OUT),
        .gtx_wait  (gtx_wait),
        .rxdv      (rxdv_snapr[5]),
        .rxcomma   (rxcomma_snapr[5]),
        .check_ok  (check_ok_snapr[5]),
        .check_bad (check_bad_snapr[5]),
        .good_byte (good_byte[5]),
        .bad_byte  (bad_byte[5]),
        .lost_byte (lost_byte[5]),
        .err_count (errcount5),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .RXCLKCORCNT_OUT                (GTX9_RXCLKCORCNT_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEREALIGN_OUT              (GTX9_RXBYTEREALIGN_OUT),
        .RXCOMMADET_OUT                 (GTX9_RXCOMMADET_OUT),
        .RXENMCOMMAALIGN_IN             (GTX9_RXENMCOMMAALIGN_IN),
        .RXENPCOMMAALIGN_IN             (GTX9_RXENPCOMMAALIGN_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA_OUT                     (),
        .RXCHARISK_OUT                  (),
        .RXRESET_IN                     (GTX9_RXRESET_IN),
        .RXUSRCLK2_IN                   (GTX9_RXUSRCLK2_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXCDRRESET_IN                  (GTX9_RXCDRRESET_IN),
        .RXN_IN                         (GTX9_RXN_IN),
        .RXP_IN                         (GTX9_RXP_IN),
        //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg        .RXBUFSTATUS_OUT                (GTX9_RXBUFSTATUS_OUT),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .RXLOSSOFSYNC_OUT               (GTX9_RXLOSSOFSYNC_OUT),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTXRXRESET_IN                  (GTX9_GTXRXRESET_IN),
        .MGTREFCLKRX_IN                 ({tied_to_ground_i , GTX9_MGTREFCLKRX_IN}),
        .PLLRXRESET_IN                  (GTX9_PLLRXRESET_IN),
        .RXPLLLKDET_OUT                 (GTX9_RXPLLLKDET_OUT),
        .RXRESETDONE_OUT                (GTX9_RXRESETDONE_OUT),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .RXVALID_OUT                    (GTX9_RXVALID_OUT),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY_IN                  (GTX9_RXPOLARITY_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .iseed                       (GTX9_SEED_IN),
        .rxseed                      (GTX9_RXSEED),
        .force_error                 (gtx9_force_error),
        .TXOUTCLK_OUT                   (GTX9_TXOUTCLK_OUT),
        .TXRESET_IN                     (GTX9_TXRESET_IN),
        .TXUSRCLK2_IN                   (GTX9_TXUSRCLK2_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .TXN_OUT                        (GTX9_TXN_OUT),
        .TXP_OUT                        (GTX9_TXP_OUT),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .TXDLYALIGNDISABLE_IN           (GTX9_TXDLYALIGNDISABLE_IN),
        .TXDLYALIGNMONENB_IN            (GTX9_TXDLYALIGNMONENB_IN),
        .TXDLYALIGNMONITOR_OUT          (GTX9_TXDLYALIGNMONITOR_OUT),
        .TXDLYALIGNRESET_IN             (GTX9_TXDLYALIGNRESET_IN),
        .TXENPMAPHASEALIGN_IN           (GTX9_TXENPMAPHASEALIGN_IN),
        .TXPMASETPHASE_IN               (GTX9_TXPMASETPHASE_IN),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTXTXRESET_IN                  (GTX9_GTXTXRESET_IN),
        .MGTREFCLKTX_IN                 ({tied_to_ground_i , GTX9_MGTREFCLKRX_IN}),
        .PLLTXRESET_IN                  (tied_to_ground_i),
        .TXPLLLKDET_OUT                 (),
        .TXRESETDONE_OUT                (GTX9_TXRESETDONE_OUT)
    );

//_________________________________________________________________________
//_________________________________________________________________________
//GTX10  (X0Y10)  TX5-fiber10 + RX6-fiber11[boardRX10]
    SNAP12_T20R20_GTX #
    (
        // Simulation attributes
        .GTX_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        // Share RX PLL parameter
        .GTX_TX_CLK_SOURCE           ("RXPLL"),
        // Save power parameter
        // old .GTX_POWER_SAVE              (10'b0000100100)
// new default        
        .GTX_POWER_SAVE              (10'b0000110000)
    )
    gtx10_snap12_t20r20_i
    (
        //---------------------- Loopback and Powerdown Ports ----------------------
        .RXPOWERDOWN_IN                 (low2),
        .TXPOWERDOWN_IN                 (low2),
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg        .RXCHARISCOMMA_OUT              (GTX10_RXCHARISCOMMA_OUT),
//jg        .RXCHARISK_OUT                  (GTX10_RXCHARISK_OUT),
//jg        .RXDISPERR_OUT                  (GTX10_RXDISPERR_OUT),
//jg        .RXNOTINTABLE_OUT               (GTX10_RXNOTINTABLE_OUT),
        .gtx_wait  (gtx_wait),
        .rxdv      (rxdv_snapr[6]),
        .rxcomma   (rxcomma_snapr[6]),
        .check_ok  (check_ok_snapr[6]),
        .check_bad (check_bad_snapr[6]),
        .good_byte (good_byte[6]),
        .bad_byte  (bad_byte[6]),
        .lost_byte (lost_byte[6]),
        .err_count (errcount6),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .RXCLKCORCNT_OUT                (GTX10_RXCLKCORCNT_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEREALIGN_OUT              (GTX10_RXBYTEREALIGN_OUT),
        .RXCOMMADET_OUT                 (GTX10_RXCOMMADET_OUT),
        .RXENMCOMMAALIGN_IN             (GTX10_RXENMCOMMAALIGN_IN),
        .RXENPCOMMAALIGN_IN             (GTX10_RXENPCOMMAALIGN_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA_OUT                     (),
        .RXCHARISK_OUT                  (),
        .RXRESET_IN                     (GTX10_RXRESET_IN),
        .RXUSRCLK2_IN                   (GTX10_RXUSRCLK2_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXCDRRESET_IN                  (GTX10_RXCDRRESET_IN),
        .RXN_IN                         (GTX10_RXN_IN),
        .RXP_IN                         (GTX10_RXP_IN),
        //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg        .RXBUFSTATUS_OUT                (GTX10_RXBUFSTATUS_OUT),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .RXLOSSOFSYNC_OUT               (GTX10_RXLOSSOFSYNC_OUT),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTXRXRESET_IN                  (GTX10_GTXRXRESET_IN),
        .MGTREFCLKRX_IN                 ({tied_to_ground_i , GTX10_MGTREFCLKRX_IN}),
        .PLLRXRESET_IN                  (GTX10_PLLRXRESET_IN),
        .RXPLLLKDET_OUT                 (GTX10_RXPLLLKDET_OUT),
        .RXRESETDONE_OUT                (GTX10_RXRESETDONE_OUT),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .RXVALID_OUT                    (GTX10_RXVALID_OUT),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY_IN                  (GTX10_RXPOLARITY_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .iseed                       (GTX10_SEED_IN),
        .rxseed                      (GTX10_RXSEED),
        .force_error                 (gtx10_force_error),
        .TXOUTCLK_OUT                   (GTX10_TXOUTCLK_OUT),
        .TXRESET_IN                     (GTX10_TXRESET_IN),
        .TXUSRCLK2_IN                   (GTX10_TXUSRCLK2_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .TXN_OUT                        (GTX10_TXN_OUT),
        .TXP_OUT                        (GTX10_TXP_OUT),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .TXDLYALIGNDISABLE_IN           (GTX10_TXDLYALIGNDISABLE_IN),
        .TXDLYALIGNMONENB_IN            (GTX10_TXDLYALIGNMONENB_IN),
        .TXDLYALIGNMONITOR_OUT          (GTX10_TXDLYALIGNMONITOR_OUT),
        .TXDLYALIGNRESET_IN             (GTX10_TXDLYALIGNRESET_IN),
        .TXENPMAPHASEALIGN_IN           (GTX10_TXENPMAPHASEALIGN_IN),
        .TXPMASETPHASE_IN               (GTX10_TXPMASETPHASE_IN),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTXTXRESET_IN                  (GTX10_GTXTXRESET_IN),
        .MGTREFCLKTX_IN                 ({tied_to_ground_i , GTX10_MGTREFCLKRX_IN}),
        .PLLTXRESET_IN                  (tied_to_ground_i),
        .TXPLLLKDET_OUT                 (),
        .TXRESETDONE_OUT                (GTX10_TXRESETDONE_OUT)
    );

//_________________________________________________________________________
//_________________________________________________________________________
//GTX11  (X0Y11)  TX6-fiber11 + RX7-fiber12[boardRX11]
    SNAP12_T20R20_GTX #
    (
        // Simulation attributes
        .GTX_SIM_GTXRESET_SPEEDUP   (WRAPPER_SIM_GTXRESET_SPEEDUP),
        // Share RX PLL parameter
        .GTX_TX_CLK_SOURCE           ("RXPLL"),
        // Save power parameter
        // old .GTX_POWER_SAVE              (10'b0000100100)
// new default       
        .GTX_POWER_SAVE              (10'b0000110000)
    )
    gtx11_snap12_t20r20_i
    (
        //---------------------- Loopback and Powerdown Ports ----------------------
        .RXPOWERDOWN_IN                 (low2),
        .TXPOWERDOWN_IN                 (low2),
        //--------------------- Receive Ports - 8b10b Decoder ----------------------
//jg        .RXCHARISCOMMA_OUT              (GTX11_RXCHARISCOMMA_OUT),
//jg        .RXCHARISK_OUT                  (GTX11_RXCHARISK_OUT),
//jg        .RXDISPERR_OUT                  (GTX11_RXDISPERR_OUT),
//jg        .RXNOTINTABLE_OUT               (GTX11_RXNOTINTABLE_OUT),
        .gtx_wait  (gtx_wait),
        .rxdv      (rxdv_snapr[7]),
        .rxcomma   (rxcomma_snapr[7]),
        .check_ok  (check_ok_snapr[7]),
        .check_bad (check_bad_snapr[7]),
        .good_byte (good_byte[7]),
        .bad_byte  (bad_byte[7]),
        .lost_byte (lost_byte[7]),
        .err_count (errcount7),
        //----------------- Receive Ports - Clock Correction Ports -----------------
        .RXCLKCORCNT_OUT                (GTX11_RXCLKCORCNT_OUT),
        //------------- Receive Ports - Comma Detection and Alignment --------------
        .RXBYTEREALIGN_OUT              (GTX11_RXBYTEREALIGN_OUT),
        .RXCOMMADET_OUT                 (GTX11_RXCOMMADET_OUT),
        .RXENMCOMMAALIGN_IN             (GTX11_RXENMCOMMAALIGN_IN),
        .RXENPCOMMAALIGN_IN             (GTX11_RXENPCOMMAALIGN_IN),
        //----------------- Receive Ports - RX Data Path interface -----------------
        .RXDATA_OUT                     (),
        .RXCHARISK_OUT                  (),
        .RXRESET_IN                     (GTX11_RXRESET_IN),
        .RXUSRCLK2_IN                   (GTX11_RXUSRCLK2_IN),
        //----- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        .RXCDRRESET_IN                  (GTX11_RXCDRRESET_IN),
        .RXN_IN                         (GTX11_RXN_IN),
        .RXP_IN                         (GTX11_RXP_IN),
        //------ Receive Ports - RX Elastic Buffer and Phase Alignment Ports -------
//jg        .RXBUFSTATUS_OUT                (GTX11_RXBUFSTATUS_OUT),
        //------------- Receive Ports - RX Loss-of-sync State Machine --------------
        .RXLOSSOFSYNC_OUT               (GTX11_RXLOSSOFSYNC_OUT),
        //---------------------- Receive Ports - RX PLL Ports ----------------------
        .GTXRXRESET_IN                  (GTX11_GTXRXRESET_IN),
        .MGTREFCLKRX_IN                 ({tied_to_ground_i , GTX11_MGTREFCLKRX_IN}),
        .PLLRXRESET_IN                  (GTX11_PLLRXRESET_IN),
        .RXPLLLKDET_OUT                 (GTX11_RXPLLLKDET_OUT),
        .RXRESETDONE_OUT                (GTX11_RXRESETDONE_OUT),
        //------------ Receive Ports - RX Pipe Control for PCI Express -------------
        .RXVALID_OUT                    (GTX11_RXVALID_OUT),
        //--------------- Receive Ports - RX Polarity Control Ports ----------------
        .RXPOLARITY_IN                  (GTX11_RXPOLARITY_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .iseed                       (GTX11_SEED_IN),
        .rxseed                      (GTX11_RXSEED),
        .force_error                 (gtx11_force_error),
        .TXOUTCLK_OUT                   (GTX11_TXOUTCLK_OUT),
        .TXRESET_IN                     (GTX11_TXRESET_IN),
        .TXUSRCLK2_IN                   (GTX11_TXUSRCLK2_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .TXN_OUT                        (GTX11_TXN_OUT),
        .TXP_OUT                        (GTX11_TXP_OUT),
        //------ Transmit Ports - TX Elastic Buffer and Phase Alignment Ports ------
        .TXDLYALIGNDISABLE_IN           (GTX11_TXDLYALIGNDISABLE_IN),
        .TXDLYALIGNMONENB_IN            (GTX11_TXDLYALIGNMONENB_IN),
        .TXDLYALIGNMONITOR_OUT          (GTX11_TXDLYALIGNMONITOR_OUT),
        .TXDLYALIGNRESET_IN             (GTX11_TXDLYALIGNRESET_IN),
        .TXENPMAPHASEALIGN_IN           (GTX11_TXENPMAPHASEALIGN_IN),
        .TXPMASETPHASE_IN               (GTX11_TXPMASETPHASE_IN),
        //--------------------- Transmit Ports - TX PLL Ports ----------------------
        .GTXTXRESET_IN                  (GTX11_GTXTXRESET_IN),
        .MGTREFCLKTX_IN                 ({tied_to_ground_i , GTX11_MGTREFCLKRX_IN}),
        .PLLTXRESET_IN                  (tied_to_ground_i),
        .TXPLLLKDET_OUT                 (),
        .TXRESETDONE_OUT                (GTX11_TXRESETDONE_OUT)
    );

endmodule
